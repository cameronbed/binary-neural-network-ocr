`ifndef SYNTHESIS
`include "Conv2d_MaxPool2d.sv"
`include "FC.sv"
`include "Comparator.sv"
`endif

module bnn_top #(
    parameter int CONV1_IMG_IN_SIZE = 30,
    parameter int CONV1_IMG_OUT_SIZE = CONV1_IMG_IN_SIZE - 2,
    parameter int POOL1_IMG_OUT_SIZE = CONV1_IMG_OUT_SIZE / 2,
    parameter int CONV2_IMG_OUT_SIZE = POOL1_IMG_OUT_SIZE - 2,
    parameter int POOL2_IMG_OUT_SIZE = CONV2_IMG_OUT_SIZE / 2,
    parameter int CONV1_IC = 1,
    parameter int CONV1_OC = 16,
    parameter int CONV2_OC = 16,
    parameter int FC_OC = 10,  // num classes
    parameter int FC_IC = POOL2_IMG_OUT_SIZE * POOL2_IMG_OUT_SIZE * CONV2_OC,
    parameter int OUTPUT_BIT = $clog2(FC_OC + 1)  // num of bits to enumerate each class
) (

    input logic [CONV1_IMG_IN_SIZE*CONV1_IMG_IN_SIZE-1:0] conv1_img_in[0:CONV1_IC-1],
    input logic clk,
    input logic data_in_ready,
    output logic [OUTPUT_BIT-1:0] result,
    output logic data_out_ready
);
  // assign conv1_img_in = img_in;
  (* rom_style = "block" *)
  logic [CONV1_IC*9-1:0] conv1_weights[0:CONV1_OC-1] = {
    9'h28,
    9'h1c4,
    9'h17d,
    9'h1e2,
    9'haf,
    9'hb1,
    9'hb5,
    9'h1ca,
    9'h1b1,
    9'h79,
    9'h6d,
    9'h1d5,
    9'h145,
    9'h158,
    9'ha0,
    9'h11c
  };
  (* rom_style = "block" *)
  logic [CONV1_OC*9-1:0] conv2_weights[0:CONV2_OC-1] = {
    144'h984335a06929ef25208409fdd624c6748e9b,
    144'h68108466d749bd0212f066503bb9ca085040,
    144'h8768853822e3d825008e080023c3e4701620,
    144'h179df335e6a6dbec6b6c87c5cab6884c9c82,
    144'h7515da842de59a4cefa267e1f5fd3949be1b,
    144'h68ae471f7e1e7e9fced5c121dabc6077c03,
    144'h942ef0d88693634c1f2d8d274c0802bb77af,
    144'h604e20512e026bb6f2d2b1831f1a97122b4e,
    144'h8f296b13a8527fff24fcba72e9b8f14780f6,
    144'h9c8edfc1d770273aee76300554bd01007901,
    144'h2e47a5db0eae65c9393c6ddc3f0c95eca80,
    144'h7d50100289b3d1364ac308060187301089bc,
    144'hf2ffd0a10994db50c104100d407520dea2f8,
    144'hba3e10666819e0c1f984803fd01ac69d02,
    144'h9eb9a03a85d5a100d42254c10277183d062,
    144'h87a21004884c742e41665be8521c90db00c3
  };
  (* rom_style = "block" *)
  logic signed [15:0] fc_weights[0:FC_IC*FC_OC-1] = {
    16'h0,
    16'hffe7,
    16'h14,
    16'h1b,
    16'hc,
    16'hf,
    16'h3,
    16'hffe6,
    16'hfffc,
    16'ha,
    16'h5,
    16'ha,
    16'h2,
    16'hfff8,
    16'h0,
    16'hffe8,
    16'h1a,
    16'hfff7,
    16'ha,
    16'hfff9,
    16'h3,
    16'h16,
    16'hfffe,
    16'hfff6,
    16'hfff8,
    16'hffed,
    16'hfff2,
    16'hfff8,
    16'h13,
    16'he,
    16'hd,
    16'h7,
    16'hfffa,
    16'hffed,
    16'h3,
    16'h16,
    16'hfff0,
    16'h15,
    16'hfff5,
    16'h15,
    16'h4,
    16'h7,
    16'hfffc,
    16'hfffc,
    16'h26,
    16'h2e,
    16'h27,
    16'hc,
    16'hfff7,
    16'h1f,
    16'hb,
    16'hffe2,
    16'h2b,
    16'h29,
    16'h1b,
    16'h18,
    16'hffd7,
    16'hffce,
    16'hfffe,
    16'hf,
    16'hfff8,
    16'h19,
    16'h1e,
    16'hffe6,
    16'hffde,
    16'h15,
    16'h1b,
    16'h15,
    16'h27,
    16'h7,
    16'hfff0,
    16'h0,
    16'hfffd,
    16'hfff6,
    16'hfff4,
    16'hfff9,
    16'hffe5,
    16'hffe1,
    16'h1,
    16'hfffc,
    16'h5,
    16'h11,
    16'hd,
    16'hffec,
    16'hffe9,
    16'hffef,
    16'h1d,
    16'hfffe,
    16'hfff0,
    16'h1,
    16'hffe6,
    16'h4,
    16'hffe7,
    16'hffe3,
    16'h33,
    16'hf,
    16'h8,
    16'h6,
    16'hfff3,
    16'h21,
    16'ha,
    16'h14,
    16'h0,
    16'h1b,
    16'hf,
    16'h7,
    16'hfff6,
    16'h4,
    16'hb,
    16'hfff9,
    16'hffe1,
    16'h1b,
    16'ha,
    16'h9,
    16'hffea,
    16'hfff0,
    16'h9,
    16'hfff9,
    16'hfff7,
    16'hfffe,
    16'hfffb,
    16'hfffa,
    16'h7,
    16'hffea,
    16'hfff0,
    16'hffc0,
    16'hfff5,
    16'hfff2,
    16'h12,
    16'hffe8,
    16'h2,
    16'h2,
    16'hfff1,
    16'hd,
    16'h15,
    16'h14,
    16'h1e,
    16'h8,
    16'h0,
    16'h18,
    16'h1b,
    16'hfffd,
    16'h1a,
    16'hfff6,
    16'hfffb,
    16'hffd7,
    16'h19,
    16'he,
    16'hffe2,
    16'hffd8,
    16'hfffd,
    16'hd,
    16'h5,
    16'hfff4,
    16'hfff4,
    16'hfffd,
    16'hffe3,
    16'h1d,
    16'hffec,
    16'hfff0,
    16'h19,
    16'h1f,
    16'hffe9,
    16'h12,
    16'hffac,
    16'h17,
    16'h13,
    16'h4,
    16'hffe8,
    16'h1e,
    16'h12,
    16'h1d,
    16'h1,
    16'h8,
    16'hffef,
    16'h4,
    16'hfff4,
    16'h0,
    16'hffe5,
    16'hfffc,
    16'hb,
    16'hffe4,
    16'hffde,
    16'hfffa,
    16'h9,
    16'hfff5,
    16'hfffc,
    16'h3,
    16'h16,
    16'h6,
    16'h14,
    16'h1e,
    16'ha,
    16'h38,
    16'hffef,
    16'hffb6,
    16'h7,
    16'he,
    16'hfff7,
    16'h18,
    16'hfffe,
    16'h17,
    16'h27,
    16'hfffa,
    16'hfff7,
    16'hfff6,
    16'h2d,
    16'hfffa,
    16'hfffb,
    16'hfff3,
    16'hc,
    16'hfff8,
    16'hfff1,
    16'hffff,
    16'h5,
    16'hffe5,
    16'he,
    16'h2,
    16'hffe7,
    16'hfff4,
    16'h8,
    16'hfffa,
    16'hfff1,
    16'h14,
    16'hffef,
    16'hffe8,
    16'hffea,
    16'hb,
    16'h6,
    16'hfff5,
    16'h10,
    16'hfffe,
    16'hffed,
    16'hfff8,
    16'hfff2,
    16'hffee,
    16'h15,
    16'h9,
    16'hffff,
    16'h14,
    16'hffe6,
    16'h5,
    16'hfff1,
    16'h25,
    16'h18,
    16'h10,
    16'hfff7,
    16'hfff8,
    16'h11,
    16'h9,
    16'hffe6,
    16'h19,
    16'h7,
    16'hfffc,
    16'hffeb,
    16'h18,
    16'h1f,
    16'hfffe,
    16'hfff1,
    16'h4,
    16'h3,
    16'hfff8,
    16'h11,
    16'h7,
    16'h8,
    16'h1,
    16'hffe3,
    16'hffd4,
    16'h3,
    16'h9,
    16'h1,
    16'h11,
    16'hffdb,
    16'hfff7,
    16'hfff3,
    16'h0,
    16'hfff6,
    16'h22,
    16'hd,
    16'ha,
    16'hffef,
    16'hffe4,
    16'h7,
    16'hfffa,
    16'hffff,
    16'hffe9,
    16'hfff0,
    16'hfffa,
    16'h19,
    16'hffe0,
    16'h11,
    16'hfff8,
    16'hffed,
    16'hffe9,
    16'h1,
    16'hd,
    16'h11,
    16'hb,
    16'he,
    16'hfff8,
    16'ha,
    16'hfff8,
    16'h22,
    16'h2,
    16'hffdc,
    16'hfffb,
    16'hffce,
    16'hffc8,
    16'hffff,
    16'ha,
    16'hffd8,
    16'hb,
    16'hffd2,
    16'hffc1,
    16'h1a,
    16'hc,
    16'hffea,
    16'h1d,
    16'hfffc,
    16'hfff0,
    16'h24,
    16'hd,
    16'hfff6,
    16'hfffa,
    16'hfff9,
    16'hffe5,
    16'h9,
    16'hfffc,
    16'h7,
    16'hffef,
    16'hfffe,
    16'h1d,
    16'h5,
    16'hffde,
    16'hffdf,
    16'hfff6,
    16'h5,
    16'hc,
    16'h3,
    16'hff95,
    16'hffcc,
    16'hfffb,
    16'hffd1,
    16'hffe7,
    16'h18,
    16'h20,
    16'hfffb,
    16'hffee,
    16'hffd7,
    16'hffd9,
    16'h1d,
    16'hfffe,
    16'hfff7,
    16'hfff8,
    16'hfffa,
    16'hffdf,
    16'hfff4,
    16'h3,
    16'h1d,
    16'h15,
    16'h16,
    16'hffee,
    16'hffe5,
    16'hffcd,
    16'hffcf,
    16'h8,
    16'h11,
    16'hffef,
    16'hffeb,
    16'hfff8,
    16'h3,
    16'hffee,
    16'h15,
    16'hffe6,
    16'h16,
    16'h24,
    16'h1f,
    16'hfffb,
    16'hf,
    16'h35,
    16'h1f,
    16'hffde,
    16'h3,
    16'h14,
    16'h10,
    16'h1f,
    16'hfff7,
    16'hffe0,
    16'hfff7,
    16'h7,
    16'hfff9,
    16'hfffa,
    16'h14,
    16'hffe8,
    16'hf,
    16'hfff8,
    16'hf,
    16'hfffe,
    16'h1,
    16'hb,
    16'h1,
    16'h0,
    16'h10,
    16'hffef,
    16'hffe7,
    16'hfff3,
    16'h5,
    16'hfff7,
    16'hffe9,
    16'hffec,
    16'hffda,
    16'h2a,
    16'h3,
    16'hffcd,
    16'hfffc,
    16'hffc3,
    16'hffdf,
    16'h1,
    16'hffef,
    16'hfffe,
    16'hfff0,
    16'hffe0,
    16'hffec,
    16'hfff6,
    16'h15,
    16'h18,
    16'he,
    16'h19,
    16'h14,
    16'hfff7,
    16'h16,
    16'h10,
    16'hfff0,
    16'he,
    16'hc,
    16'h5,
    16'hfff4,
    16'hfff6,
    16'hfff9,
    16'hfffe,
    16'hffed,
    16'hfff6,
    16'hffd3,
    16'hfff3,
    16'hd,
    16'hffff,
    16'hfff7,
    16'h18,
    16'hffed,
    16'hffe1,
    16'hffea,
    16'hfff6,
    16'hffdf,
    16'h6,
    16'h6,
    16'hfffd,
    16'h7,
    16'hffec,
    16'hfff9,
    16'h3,
    16'h9,
    16'hf,
    16'hffef,
    16'h5,
    16'hffed,
    16'h0,
    16'hffea,
    16'hffea,
    16'hfff6,
    16'hffed,
    16'h8,
    16'h12,
    16'he,
    16'hc,
    16'hfff0,
    16'h1,
    16'h2e,
    16'h9,
    16'h1c,
    16'h8,
    16'hffed,
    16'h19,
    16'h2f,
    16'hffe6,
    16'h1f,
    16'h3a,
    16'hffea,
    16'h35,
    16'h21,
    16'hffca,
    16'h18,
    16'h35,
    16'he,
    16'h16,
    16'h7,
    16'hffd3,
    16'hffee,
    16'hfff6,
    16'h11,
    16'hb,
    16'hfff2,
    16'hfff6,
    16'hffe6,
    16'hfff6,
    16'h16,
    16'h10,
    16'hffff,
    16'h1f,
    16'h4,
    16'h17,
    16'hfff8,
    16'he,
    16'hb,
    16'hfff1,
    16'hfff3,
    16'hffea,
    16'hfff8,
    16'hffe5,
    16'hffeb,
    16'h29,
    16'h6,
    16'hffdf,
    16'h1,
    16'hffd6,
    16'hffe6,
    16'h19,
    16'hfff4,
    16'hffd7,
    16'h6,
    16'hfffc,
    16'hffd9,
    16'h0,
    16'h6,
    16'h1,
    16'h17,
    16'hffec,
    16'hfffc,
    16'h3,
    16'h0,
    16'hffef,
    16'h8,
    16'h13,
    16'h9,
    16'hfff3,
    16'h8,
    16'ha,
    16'h4,
    16'hfff9,
    16'hfff9,
    16'h1e,
    16'h6,
    16'hfff1,
    16'hfff1,
    16'hffff,
    16'hffdb,
    16'hfffb,
    16'h21,
    16'hfff3,
    16'hfffe,
    16'h2,
    16'hffa9,
    16'hffb0,
    16'hffdf,
    16'hffec,
    16'h12,
    16'h16,
    16'hffd8,
    16'hffca,
    16'hc,
    16'h16,
    16'h25,
    16'h22,
    16'h26,
    16'h2b,
    16'hffe3,
    16'hfff4,
    16'hfff7,
    16'hfffe,
    16'h18,
    16'h17,
    16'hffff,
    16'hfff5,
    16'hfffb,
    16'hd,
    16'h17,
    16'h29,
    16'h5,
    16'h15,
    16'h10,
    16'hfffb,
    16'hffeb,
    16'ha,
    16'hfff9,
    16'h18,
    16'hf,
    16'h6,
    16'hfffc,
    16'hd,
    16'hfffc,
    16'hffee,
    16'hfff8,
    16'h15,
    16'hffef,
    16'hf,
    16'hfff7,
    16'hffed,
    16'h8,
    16'hfffa,
    16'h0,
    16'h1a,
    16'hb,
    16'h14,
    16'hfff6,
    16'h6,
    16'hffee,
    16'hf,
    16'hffff,
    16'hfff0,
    16'hfff4,
    16'h7,
    16'h46,
    16'h1a,
    16'hfff5,
    16'hffee,
    16'hfff1,
    16'hffe2,
    16'h2,
    16'h1c,
    16'hfff9,
    16'hffe4,
    16'h9,
    16'hffec,
    16'hfffe,
    16'hfff6,
    16'hfff4,
    16'h8,
    16'hfff5,
    16'hfff3,
    16'h0,
    16'h1b,
    16'hfffc,
    16'h3,
    16'hffe6,
    16'h2,
    16'he,
    16'h16,
    16'h9,
    16'hfff0,
    16'ha,
    16'hfff2,
    16'hfff8,
    16'h17,
    16'h12,
    16'h2d,
    16'hc,
    16'hfff8,
    16'hfff4,
    16'hfffe,
    16'h9,
    16'hfff6,
    16'hb,
    16'hffea,
    16'hfff2,
    16'h9,
    16'hffef,
    16'hffec,
    16'h13,
    16'hffc7,
    16'h21,
    16'h17,
    16'hffd8,
    16'hfff9,
    16'hffdb,
    16'hffe1,
    16'h20,
    16'hffc0,
    16'h5,
    16'h21,
    16'hf,
    16'hffff,
    16'hfffe,
    16'hffef,
    16'h13,
    16'hfff5,
    16'hf,
    16'hfff4,
    16'hfffd,
    16'hffd9,
    16'hfff6,
    16'h4,
    16'h1,
    16'hffed,
    16'hffb8,
    16'h16,
    16'hffdc,
    16'hfffb,
    16'h0,
    16'h7,
    16'h3,
    16'h6,
    16'hffe8,
    16'hffd7,
    16'he,
    16'hffe7,
    16'hffe9,
    16'hfff6,
    16'hfffd,
    16'hfff5,
    16'hfffc,
    16'hffe2,
    16'hffed,
    16'hffff,
    16'hffe9,
    16'h11,
    16'h1f,
    16'h0,
    16'ha,
    16'hffdf,
    16'hfff8,
    16'h25,
    16'hfff7,
    16'hffe9,
    16'hffd4,
    16'hfffc,
    16'h4,
    16'hffe1,
    16'hfff6,
    16'hffaf,
    16'hfff1,
    16'hffca,
    16'hffdf,
    16'hffff,
    16'hc,
    16'hffe3,
    16'h1c,
    16'hffeb,
    16'hffbd,
    16'hffe7,
    16'hfff8,
    16'hffe8,
    16'h4,
    16'hffc5,
    16'hffd4,
    16'h6,
    16'h9,
    16'hffef,
    16'hffe9,
    16'hffd0,
    16'h6,
    16'hfff9,
    16'ha,
    16'hffe3,
    16'hffef,
    16'hffe3,
    16'h9,
    16'h1,
    16'hfffa,
    16'hfff4,
    16'hffd9,
    16'h7,
    16'hfffd,
    16'h1,
    16'h0,
    16'hffe1,
    16'hffd6,
    16'h7,
    16'hffc8,
    16'hffe1,
    16'hfff1,
    16'hffc8,
    16'hfff8,
    16'h4,
    16'hffc6,
    16'hffe7,
    16'hffee,
    16'hffcb,
    16'hfffc,
    16'h6,
    16'hffc3,
    16'hfffd,
    16'h2,
    16'ha,
    16'hffef,
    16'hffcf,
    16'h17,
    16'h0,
    16'hf,
    16'hffe3,
    16'hffde,
    16'hffc2,
    16'hffe4,
    16'h0,
    16'h1a,
    16'h10,
    16'h7,
    16'hfff5,
    16'hffee,
    16'hfff6,
    16'hfff7,
    16'hffeb,
    16'hfffe,
    16'hf,
    16'h10,
    16'h0,
    16'hf,
    16'h1,
    16'ha,
    16'hf,
    16'ha,
    16'h1a,
    16'h4,
    16'h0,
    16'hfff3,
    16'h8,
    16'hfff2,
    16'h15,
    16'h0,
    16'h14,
    16'h1,
    16'hffed,
    16'hfff8,
    16'h13,
    16'h9,
    16'hc,
    16'hfff5,
    16'hf,
    16'hfff7,
    16'h3,
    16'hfff0,
    16'hffef,
    16'hffd1,
    16'hffdb,
    16'hfff2,
    16'hffee,
    16'h6,
    16'hfff9,
    16'hfff8,
    16'h1a,
    16'hffd0,
    16'hffdf,
    16'hffee,
    16'hffd8,
    16'hfffe,
    16'h13,
    16'hffcd,
    16'h5,
    16'hffdd,
    16'hffeb,
    16'h11,
    16'hffdd,
    16'hffdb,
    16'h0,
    16'h4,
    16'hfff0,
    16'h2,
    16'h7,
    16'h29,
    16'hfffa,
    16'hfffb,
    16'hfff3,
    16'hfff0,
    16'hffef,
    16'hfffe,
    16'hfff0,
    16'hffeb,
    16'hffeb,
    16'hffee,
    16'hfffe,
    16'h11,
    16'h2,
    16'h16,
    16'hfff7,
    16'hfff5,
    16'hffc4,
    16'hffe5,
    16'hffe4,
    16'hb,
    16'hfffe,
    16'hffd6,
    16'h11,
    16'hffee,
    16'hffef,
    16'he,
    16'h18,
    16'hffb8,
    16'h7,
    16'hffee,
    16'hfff2,
    16'h11,
    16'hfff4,
    16'hffc7,
    16'hfff8,
    16'hb,
    16'hd,
    16'hfffd,
    16'hb,
    16'hfff3,
    16'hfff6,
    16'hffe6,
    16'h13,
    16'h7,
    16'h11,
    16'hc,
    16'hfff1,
    16'hfff8,
    16'h16,
    16'hfff7,
    16'hffe5,
    16'hfff3,
    16'h11,
    16'ha,
    16'hfff6,
    16'h1c,
    16'h10,
    16'hffe1,
    16'hfff5,
    16'h5,
    16'h7,
    16'hfffb,
    16'ha,
    16'hffdb,
    16'hfff8,
    16'hfffa,
    16'h1a,
    16'hfffa,
    16'h29,
    16'hffe8,
    16'hd,
    16'hfffa,
    16'h5,
    16'h3,
    16'hffde,
    16'h1,
    16'hffdd,
    16'hffef,
    16'h1,
    16'h16,
    16'h3,
    16'hd,
    16'he,
    16'h9,
    16'hffef,
    16'hfff0,
    16'hfffd,
    16'h0,
    16'hffd3,
    16'hfff6,
    16'hfff8,
    16'hfff7,
    16'h12,
    16'hffcc,
    16'hc,
    16'hfff6,
    16'hc,
    16'hb,
    16'hfffa,
    16'h8,
    16'h2,
    16'hffed,
    16'hffe3,
    16'h5,
    16'h1,
    16'h5,
    16'h1,
    16'hfff7,
    16'hc,
    16'h1f,
    16'h11,
    16'h0,
    16'hffe2,
    16'hfffe,
    16'h1a,
    16'h16,
    16'h2,
    16'hfff5,
    16'hfffe,
    16'hffed,
    16'hffea,
    16'hd,
    16'hfffe,
    16'h1,
    16'hfffc,
    16'hffea,
    16'h9,
    16'hfff3,
    16'h10,
    16'h15,
    16'h1,
    16'h18,
    16'hfff9,
    16'h9,
    16'hc,
    16'hfff8,
    16'h5,
    16'h18,
    16'hfffa,
    16'h2,
    16'hffe6,
    16'hfff2,
    16'h21,
    16'h3,
    16'hfff7,
    16'hfff6,
    16'h16,
    16'h17,
    16'h27,
    16'h4,
    16'h19,
    16'hd,
    16'h1,
    16'h14,
    16'h1,
    16'h3,
    16'h1b,
    16'hfff7,
    16'h1d,
    16'hfff0,
    16'hffed,
    16'hffda,
    16'h15,
    16'hfff9,
    16'h11,
    16'hfff0,
    16'hffe9,
    16'h8,
    16'hfff6,
    16'h8,
    16'h6,
    16'hfffa,
    16'h12,
    16'hfff2,
    16'hfff1,
    16'h12,
    16'hfff2,
    16'h5,
    16'hfffc,
    16'hfff0,
    16'hffef,
    16'h4,
    16'hfff1,
    16'hfff6,
    16'hfff6,
    16'h10,
    16'h7,
    16'hffe6,
    16'hffe8,
    16'h25,
    16'h4a,
    16'h13,
    16'he,
    16'h2,
    16'hffe9,
    16'h2b,
    16'h5d,
    16'h2,
    16'h16,
    16'hfffa,
    16'h10,
    16'hffe8,
    16'h34,
    16'hd,
    16'hfff0,
    16'ha,
    16'hffe3,
    16'h12,
    16'h28,
    16'hffe6,
    16'hfff0,
    16'hffee,
    16'h1e,
    16'h28,
    16'he,
    16'hffdb,
    16'hfff6,
    16'h17,
    16'hffef,
    16'h7,
    16'hffeb,
    16'h7,
    16'hfffc,
    16'h4,
    16'h8,
    16'hfff0,
    16'hc,
    16'h5,
    16'hfffd,
    16'hfffe,
    16'hc,
    16'h24,
    16'h1e,
    16'hffd9,
    16'hfff3,
    16'h7,
    16'h1,
    16'h36,
    16'hffd9,
    16'h0,
    16'hfffa,
    16'hfffa,
    16'hc,
    16'h2d,
    16'hfff2,
    16'h7,
    16'hfff0,
    16'hffed,
    16'h3,
    16'h1d,
    16'h16,
    16'hffd8,
    16'hd,
    16'h1,
    16'hfff6,
    16'h19,
    16'h6,
    16'hffff,
    16'hfff9,
    16'h0,
    16'hfff3,
    16'h3,
    16'h5,
    16'hffec,
    16'h9,
    16'hffff,
    16'hfffd,
    16'hffff,
    16'hffdd,
    16'h4,
    16'hb,
    16'h0,
    16'h2,
    16'h1a,
    16'hfffc,
    16'hffe8,
    16'hffe2,
    16'h0,
    16'hffe4,
    16'h15,
    16'hfff6,
    16'hffe5,
    16'h8,
    16'hfff1,
    16'hfff7,
    16'h14,
    16'h11,
    16'hfff5,
    16'hb,
    16'h9,
    16'h19,
    16'hfffc,
    16'hfffe,
    16'h1f,
    16'hffff,
    16'hc,
    16'hffed,
    16'hffef,
    16'h8,
    16'hfffa,
    16'h9,
    16'h8,
    16'h5,
    16'h13,
    16'hfffa,
    16'hb,
    16'h4,
    16'hfff1,
    16'h14,
    16'h3,
    16'hfffe,
    16'hfffb,
    16'hf,
    16'hfffd,
    16'h2,
    16'hfff7,
    16'h0,
    16'h8,
    16'h8,
    16'h13,
    16'hffdf,
    16'hffeb,
    16'he,
    16'h10,
    16'h18,
    16'hfff9,
    16'hf,
    16'hffeb,
    16'h10,
    16'h7,
    16'hfff1,
    16'h17,
    16'h7,
    16'h15,
    16'h17,
    16'hffee,
    16'hfffb,
    16'hfffc,
    16'hffeb,
    16'he,
    16'h22,
    16'h30,
    16'hfffc,
    16'hffff,
    16'hffd5,
    16'hffd1,
    16'hffe8,
    16'hfffd,
    16'hfff7,
    16'hfff5,
    16'hffed,
    16'hffe4,
    16'hfff8,
    16'hffd4,
    16'hffec,
    16'h21,
    16'h21,
    16'h32,
    16'h11,
    16'hffec,
    16'h9,
    16'h3,
    16'hfffa,
    16'h10,
    16'he,
    16'hfff7,
    16'hfff1,
    16'h14,
    16'hfffb,
    16'ha,
    16'hffe8,
    16'hffd7,
    16'hffe4,
    16'h5,
    16'hf,
    16'h28,
    16'ha,
    16'hffe1,
    16'hffe4,
    16'h14,
    16'hfffb,
    16'hffe6,
    16'hfffc,
    16'hfff5,
    16'hffff,
    16'hffd5,
    16'hffe6,
    16'he,
    16'h19,
    16'h17,
    16'h21,
    16'h4,
    16'hfff2,
    16'he,
    16'hfff0,
    16'h4,
    16'h35,
    16'h26,
    16'h9,
    16'hffca,
    16'hfff9,
    16'hfff9,
    16'h19,
    16'hfff6,
    16'h7,
    16'hfff4,
    16'h22,
    16'h6,
    16'hffee,
    16'h1c,
    16'ha,
    16'h7,
    16'h14,
    16'hffd5,
    16'hffcc,
    16'h14,
    16'h17,
    16'hfffe,
    16'hb,
    16'hffe4,
    16'hffe5,
    16'h3,
    16'hfff0,
    16'hfff7,
    16'h9,
    16'he,
    16'h39,
    16'h1,
    16'hfffd,
    16'hffef,
    16'hfffb,
    16'h38,
    16'h4c,
    16'hb,
    16'h16,
    16'hffef,
    16'hffd5,
    16'h13,
    16'h1b,
    16'h5,
    16'h11,
    16'h1f,
    16'hffdd,
    16'hffef,
    16'hffd7,
    16'h9,
    16'hfffe,
    16'h26,
    16'hffea,
    16'hffde,
    16'hfff5,
    16'h1c,
    16'hfff6,
    16'he,
    16'hfffc,
    16'hffec,
    16'h7,
    16'h5,
    16'h8,
    16'h19,
    16'hfffb,
    16'ha,
    16'h2a,
    16'hfff5,
    16'h10,
    16'hfff3,
    16'h3f,
    16'h35,
    16'h49,
    16'hf,
    16'h5,
    16'h3,
    16'h16,
    16'h29,
    16'h2a,
    16'hd,
    16'hffff,
    16'h13,
    16'hffd3,
    16'hffee,
    16'h9,
    16'hfff0,
    16'hfff2,
    16'hffb7,
    16'h2,
    16'hffff,
    16'hfff6,
    16'hfffe,
    16'hffff,
    16'hffe6,
    16'h16,
    16'hfffd,
    16'hfff3,
    16'h22,
    16'ha,
    16'h2b,
    16'h17,
    16'hfff2,
    16'hffff,
    16'hffff,
    16'hf,
    16'hfff9,
    16'hffe6,
    16'h1b,
    16'h1b,
    16'h3,
    16'hffe3,
    16'hffe0,
    16'hffe6,
    16'hfff1,
    16'hffee,
    16'h1b,
    16'hfffc,
    16'h15,
    16'h1,
    16'h17,
    16'hffea,
    16'h13,
    16'hfff9,
    16'hfffb,
    16'hffd3,
    16'hffe8,
    16'h12,
    16'hffea,
    16'h6,
    16'hfffc,
    16'h1c,
    16'hfffe,
    16'hfff9,
    16'h0,
    16'hfff6,
    16'hffeb,
    16'hffff,
    16'h2,
    16'hfffa,
    16'h1,
    16'h1a,
    16'h7,
    16'hffe7,
    16'hfffa,
    16'h6,
    16'hfff3,
    16'h2,
    16'hfff5,
    16'hfff4,
    16'h8,
    16'hfff4,
    16'hfffa,
    16'hfff0,
    16'hb,
    16'h11,
    16'h2,
    16'hffe6,
    16'hfff0,
    16'hfff7,
    16'hffff,
    16'h4,
    16'h14,
    16'hffd5,
    16'hfffe,
    16'h4,
    16'h23,
    16'h10,
    16'hffdf,
    16'hfff5,
    16'h4,
    16'hffed,
    16'hffff,
    16'h12,
    16'hffe6,
    16'h13,
    16'h18,
    16'h7,
    16'hfffa,
    16'hc,
    16'h44,
    16'h37,
    16'h13,
    16'hfff9,
    16'hfff8,
    16'h0,
    16'hd,
    16'hfff6,
    16'hffd4,
    16'h0,
    16'hfffc,
    16'hfff7,
    16'hffdd,
    16'hfff1,
    16'h6,
    16'h4,
    16'h19,
    16'h19,
    16'h1,
    16'hffed,
    16'h4a,
    16'h50,
    16'h33,
    16'h4,
    16'hffec,
    16'hd,
    16'hfffd,
    16'h11,
    16'h6,
    16'hfff4,
    16'hfff5,
    16'h5,
    16'hffe5,
    16'hffd2,
    16'hffe6,
    16'he,
    16'h17,
    16'h26,
    16'ha,
    16'h6,
    16'h6,
    16'h0,
    16'hfff8,
    16'h1e,
    16'hfff3,
    16'hfffa,
    16'hffe9,
    16'hffe2,
    16'h7,
    16'hfff1,
    16'h21,
    16'hfff0,
    16'hffd7,
    16'hffcb,
    16'hfff4,
    16'h4,
    16'h17,
    16'hfffb,
    16'h8,
    16'h25,
    16'h7,
    16'h1f,
    16'h38,
    16'h20,
    16'h12,
    16'h25,
    16'h12,
    16'hfff9,
    16'hffe9,
    16'h10,
    16'hfffd,
    16'hffe9,
    16'hffeb,
    16'hfff6,
    16'hffea,
    16'hfffd,
    16'h33,
    16'h14,
    16'h3,
    16'hfffe,
    16'hffed,
    16'h20,
    16'h14,
    16'hffe9,
    16'hffdd,
    16'h7,
    16'h8,
    16'hffff,
    16'h8,
    16'hfff7,
    16'h2,
    16'h0,
    16'h12,
    16'hfff7,
    16'hffcf,
    16'h3,
    16'h3,
    16'h5,
    16'hfffc,
    16'hffeb,
    16'hffd4,
    16'h5,
    16'h8,
    16'hffef,
    16'h0,
    16'h12,
    16'h15,
    16'h5,
    16'hffc1,
    16'hffe2,
    16'h13,
    16'h20,
    16'h2,
    16'hffeb,
    16'h0,
    16'ha,
    16'hfffc,
    16'hfffe,
    16'hf,
    16'hffff,
    16'h0,
    16'hfff8,
    16'h13,
    16'h20,
    16'h1f,
    16'ha,
    16'hfffe,
    16'hffea,
    16'h4,
    16'h55,
    16'h38,
    16'h9,
    16'hfff0,
    16'hfffe,
    16'hffef,
    16'hffd7,
    16'hffdc,
    16'hffcb,
    16'h27,
    16'h3,
    16'hffe4,
    16'hffe2,
    16'h4,
    16'hfff5,
    16'h1c,
    16'h22,
    16'h1,
    16'h2,
    16'h16,
    16'h17,
    16'h1d,
    16'he,
    16'hf,
    16'h18,
    16'hfff1,
    16'hc,
    16'hfff0,
    16'h7,
    16'hd,
    16'h1a,
    16'he,
    16'h1e,
    16'hffe3,
    16'hb,
    16'hfff1,
    16'h18,
    16'h31,
    16'hd,
    16'hfffd,
    16'h6,
    16'h5,
    16'hffd9,
    16'hffc2,
    16'hffd9,
    16'h6,
    16'h14,
    16'h1b,
    16'hfff8,
    16'hfff2,
    16'hfffb,
    16'he,
    16'h1b,
    16'hf,
    16'h1b,
    16'he,
    16'h14,
    16'hfff2,
    16'hb,
    16'hf,
    16'hfff0,
    16'hffff,
    16'hfff5,
    16'hfffa,
    16'hfff7,
    16'hfff3,
    16'hffd8,
    16'hffda,
    16'hffe8,
    16'h24,
    16'h32,
    16'hfffe,
    16'hffb0,
    16'hffc9,
    16'hffe7,
    16'h20,
    16'h16,
    16'hfff8,
    16'hfff2,
    16'h10,
    16'he,
    16'hffdf,
    16'hffb9,
    16'h15,
    16'h14,
    16'h9,
    16'hffc9,
    16'hffce,
    16'hffc8,
    16'h18,
    16'h18,
    16'hfff7,
    16'hffd9,
    16'hfffe,
    16'hc,
    16'h1,
    16'h4,
    16'h5,
    16'hffe5,
    16'hfff3,
    16'h11,
    16'hfffe,
    16'hd,
    16'ha,
    16'hd,
    16'h2,
    16'h8,
    16'h15,
    16'h34,
    16'h24,
    16'h3b,
    16'hffe6,
    16'hfffd,
    16'h13,
    16'hfff4,
    16'hffd1,
    16'hffc5,
    16'hfff4,
    16'ha,
    16'hfff9,
    16'hfffa,
    16'hffee,
    16'hfff3,
    16'h24,
    16'h22,
    16'h12,
    16'h1c,
    16'h1a,
    16'h2d,
    16'h1,
    16'h15,
    16'hfff9,
    16'h13,
    16'hd,
    16'h12,
    16'hffeb,
    16'hffee,
    16'hfff1,
    16'h24,
    16'h1b,
    16'h26,
    16'ha,
    16'hfff3,
    16'hffec,
    16'hfffe,
    16'h8,
    16'h0,
    16'hffde,
    16'hfff2,
    16'hffea,
    16'hffed,
    16'hffee,
    16'hffe4,
    16'hffe8,
    16'he,
    16'hfffe,
    16'hfffc,
    16'h5,
    16'h19,
    16'h26,
    16'h55,
    16'h0,
    16'h10,
    16'h1c,
    16'h2,
    16'h12,
    16'h25,
    16'h14,
    16'hffe7,
    16'hffec,
    16'hfff6,
    16'h6,
    16'hfff2,
    16'hd,
    16'h7,
    16'h1c,
    16'hfff4,
    16'h3,
    16'hffe9,
    16'hb,
    16'h4,
    16'hfff9,
    16'hfff7,
    16'hffea,
    16'h16,
    16'h8,
    16'ha,
    16'h14,
    16'h6,
    16'hfff7,
    16'h8,
    16'hfff9,
    16'hfffe,
    16'hfffb,
    16'hfff5,
    16'hffe5,
    16'ha,
    16'hffef,
    16'h7,
    16'h2,
    16'he,
    16'hfffc,
    16'hffe9,
    16'h11,
    16'hfffc,
    16'h7,
    16'h23,
    16'h1,
    16'h15,
    16'hfff6,
    16'hffef,
    16'hb,
    16'h27,
    16'h1a,
    16'hfff7,
    16'h10,
    16'hffb7,
    16'hffde,
    16'h1,
    16'h1,
    16'hfff5,
    16'h12,
    16'hffd3,
    16'h4,
    16'h7,
    16'h2,
    16'hfff6,
    16'h13,
    16'hfff8,
    16'hffef,
    16'hfff5,
    16'h12,
    16'hffe6,
    16'h1a,
    16'hffe7,
    16'h3,
    16'hffec,
    16'hfff9,
    16'hfffa,
    16'hffef,
    16'hc,
    16'h12,
    16'hfff3,
    16'h2,
    16'hfff7,
    16'h10,
    16'h30,
    16'hb,
    16'h2,
    16'hfffe,
    16'hfff5,
    16'h17,
    16'hffeb,
    16'hfffe,
    16'h27,
    16'h1a,
    16'hffe3,
    16'hfffc,
    16'h6,
    16'h4,
    16'hffed,
    16'hffe0,
    16'h1,
    16'h0,
    16'h8,
    16'hfff7,
    16'h11,
    16'h18,
    16'hffeb,
    16'h1a,
    16'hfff7,
    16'hffe9,
    16'hc,
    16'h0,
    16'hffee,
    16'h16,
    16'h8,
    16'hfff3,
    16'hfff7,
    16'hfffd,
    16'hffea,
    16'h36,
    16'he,
    16'hffe2,
    16'h1,
    16'hffec,
    16'hffe7,
    16'h3a,
    16'h5,
    16'hffef,
    16'h6,
    16'h25,
    16'h2d,
    16'hd,
    16'h13,
    16'hfff1,
    16'h4,
    16'h16,
    16'hffea,
    16'h8,
    16'h4,
    16'h8,
    16'h1a,
    16'hd,
    16'hffd5,
    16'h13,
    16'h25,
    16'h11,
    16'hfffc,
    16'h3c,
    16'hfffa,
    16'h19,
    16'h2a,
    16'h17,
    16'hfff7,
    16'hffee,
    16'hffe8,
    16'h31,
    16'hfff0,
    16'hd,
    16'hffe8,
    16'hffcc,
    16'hfff6,
    16'hb,
    16'hfff9,
    16'h7,
    16'ha,
    16'hffeb,
    16'hffc4,
    16'h14,
    16'hfff4,
    16'h17,
    16'hd,
    16'ha,
    16'hfff0,
    16'he,
    16'h1d,
    16'h9,
    16'h39,
    16'hffef,
    16'hffe5,
    16'h2d,
    16'h2a,
    16'h6,
    16'h5,
    16'hffe7,
    16'hffea,
    16'h1c,
    16'h8,
    16'h26,
    16'hfffc,
    16'hffe8,
    16'h0,
    16'h17,
    16'hfff3,
    16'h5,
    16'h1f,
    16'h4,
    16'hfff3,
    16'hfffe,
    16'hffd1,
    16'h13,
    16'h20,
    16'hfffb,
    16'hffde,
    16'h29,
    16'hffd8,
    16'h3,
    16'hb,
    16'h32,
    16'hfff3,
    16'h2a,
    16'h23,
    16'h14,
    16'h22,
    16'he,
    16'hfff2,
    16'h1b,
    16'h3a,
    16'h36,
    16'h27,
    16'h18,
    16'hfff1,
    16'hfffa,
    16'hfff9,
    16'h6,
    16'h4,
    16'hfff5,
    16'h15,
    16'hffed,
    16'hffec,
    16'hffdd,
    16'hffea,
    16'h6,
    16'h1,
    16'h0,
    16'hfff3,
    16'hfff7,
    16'hfffe,
    16'h10,
    16'h10,
    16'hffef,
    16'hfff2,
    16'h1d,
    16'hffe8,
    16'he,
    16'h5,
    16'hffea,
    16'hffff,
    16'hffff,
    16'hfff5,
    16'h0,
    16'h4,
    16'h5,
    16'hb,
    16'hffe6,
    16'hffef,
    16'hb,
    16'h9,
    16'h17,
    16'h7,
    16'h1e,
    16'h15,
    16'h9,
    16'hfff4,
    16'h16,
    16'hfff7,
    16'hf,
    16'h29,
    16'hffef,
    16'hffde,
    16'h2,
    16'hffdf,
    16'h9,
    16'h8,
    16'hd,
    16'h2,
    16'hfffe,
    16'h3,
    16'h19,
    16'h10,
    16'h1d,
    16'hfff5,
    16'h1e,
    16'hd,
    16'hfff9,
    16'hb,
    16'hfff4,
    16'hffe1,
    16'ha,
    16'hf,
    16'h1b,
    16'hfffb,
    16'hfffa,
    16'h2,
    16'hffe9,
    16'hfff1,
    16'hfffc,
    16'h9,
    16'hffe7,
    16'hfff7,
    16'h13,
    16'h23,
    16'h2c,
    16'h14,
    16'h9,
    16'hffed,
    16'h1f,
    16'h37,
    16'hffe1,
    16'he,
    16'hfffb,
    16'hfffe,
    16'h9,
    16'h5,
    16'hffe3,
    16'hb,
    16'hfffe,
    16'hfffe,
    16'h1,
    16'h2e,
    16'h2f,
    16'h18,
    16'h16,
    16'hffe8,
    16'hd,
    16'h19,
    16'h2b,
    16'h22,
    16'h1e,
    16'hfff2,
    16'h16,
    16'h6,
    16'hfffb,
    16'ha,
    16'h15,
    16'hfff3,
    16'hc,
    16'hfff4,
    16'h0,
    16'hfff8,
    16'h12,
    16'hfff4,
    16'ha,
    16'h23,
    16'h2e,
    16'h8,
    16'hffff,
    16'h16,
    16'h2d,
    16'h17,
    16'hffeb,
    16'hfffd,
    16'h7,
    16'hfff7,
    16'he,
    16'h2d,
    16'h43,
    16'h12,
    16'hfffa,
    16'hffee,
    16'hffff,
    16'h9,
    16'h29,
    16'h1d,
    16'h19,
    16'h10,
    16'hfff0,
    16'hfff6,
    16'h15,
    16'hfffd,
    16'hffee,
    16'h7,
    16'h2,
    16'h2f,
    16'h1f,
    16'h1a,
    16'hffef,
    16'he,
    16'ha,
    16'hd,
    16'hffdd,
    16'h16,
    16'hfff6,
    16'hfffa,
    16'hffef,
    16'hfffa,
    16'h29,
    16'h19,
    16'hc,
    16'hc,
    16'hfffa,
    16'hfff4,
    16'hffe0,
    16'h4,
    16'h8,
    16'hd,
    16'hc,
    16'h18,
    16'h2,
    16'hfff2,
    16'h20,
    16'hffe6,
    16'hfff6,
    16'hfff0,
    16'h12,
    16'h7,
    16'hb,
    16'h0,
    16'hfffd,
    16'h36,
    16'h2c,
    16'hffe3,
    16'hfff0,
    16'hffe9,
    16'h3,
    16'h47,
    16'h21,
    16'hfff9,
    16'h16,
    16'h1b,
    16'hb,
    16'h50,
    16'h4b,
    16'h23,
    16'hffea,
    16'hfff1,
    16'h0,
    16'h24,
    16'h26,
    16'hffe7,
    16'hffef,
    16'hffef,
    16'h4,
    16'hfffb,
    16'hfff1,
    16'hfff2,
    16'h9,
    16'h2,
    16'hffe7,
    16'h11,
    16'h16,
    16'h7,
    16'h9,
    16'h10,
    16'hfff2,
    16'hfff7,
    16'h11,
    16'hfff9,
    16'hffbf,
    16'hfffa,
    16'hfff2,
    16'h2c,
    16'h21,
    16'hffec,
    16'h4,
    16'h20,
    16'hfffe,
    16'hf,
    16'h1b,
    16'hb,
    16'hfff0,
    16'hffdf,
    16'hfff2,
    16'hc,
    16'h4,
    16'h0,
    16'hffef,
    16'hfff2,
    16'h13,
    16'hf,
    16'h5,
    16'hfff3,
    16'h5,
    16'hfffe,
    16'hffe7,
    16'h5,
    16'h4,
    16'h13,
    16'h9,
    16'ha,
    16'h14,
    16'hffda,
    16'hffcc,
    16'h1b,
    16'h31,
    16'h2b,
    16'h12,
    16'hffcc,
    16'hffd9,
    16'hfff4,
    16'hffeb,
    16'hffe1,
    16'h8,
    16'hfff2,
    16'hffc9,
    16'hffcf,
    16'h2,
    16'h15,
    16'hfffd,
    16'hffee,
    16'hffe4,
    16'hfff1,
    16'h1c,
    16'h14,
    16'hfffd,
    16'hfffd,
    16'hfffc,
    16'hfff6,
    16'hfff9,
    16'h0,
    16'hffed,
    16'hffe8,
    16'hfffd,
    16'hfff5,
    16'hfff1,
    16'h15,
    16'hc,
    16'hffe8,
    16'hfffc,
    16'hffd5,
    16'hffc0,
    16'hffe1,
    16'h6,
    16'h35,
    16'hf,
    16'hffc8,
    16'hc,
    16'h23,
    16'h5,
    16'h34,
    16'h28,
    16'h18,
    16'h1d,
    16'h2,
    16'hffe7,
    16'h13,
    16'h15,
    16'hffec,
    16'hfff4,
    16'hfff1,
    16'hffee,
    16'hfffb,
    16'hffe3,
    16'hffec,
    16'hd,
    16'hf,
    16'hfff3,
    16'hfffa,
    16'h12,
    16'hd,
    16'hfff4,
    16'hd,
    16'hfff8,
    16'h17,
    16'h35,
    16'hf,
    16'hffed,
    16'hfff7,
    16'hfff6,
    16'hffe4,
    16'h18,
    16'hfffc,
    16'h3,
    16'hffed,
    16'hffe8,
    16'hffe0,
    16'h2e,
    16'h2a,
    16'he,
    16'hfff7,
    16'h13,
    16'h5,
    16'h22,
    16'h6,
    16'hfffc,
    16'hffe9,
    16'h39,
    16'h12,
    16'hfff0,
    16'h2,
    16'hfff5,
    16'hffee,
    16'h10,
    16'hfff6,
    16'h7,
    16'hc,
    16'hfffe,
    16'hffeb,
    16'hffef,
    16'h5,
    16'hc,
    16'h28,
    16'hfff3,
    16'hffe1,
    16'h18,
    16'h8,
    16'hffef,
    16'h11,
    16'hf,
    16'hffeb,
    16'hfff0,
    16'hf,
    16'h14,
    16'h19,
    16'hfff2,
    16'h14,
    16'hfff4,
    16'h7,
    16'hffe8,
    16'h6,
    16'h9,
    16'h4,
    16'hffee,
    16'h7,
    16'h12,
    16'hfffc,
    16'hfff4,
    16'hffeb,
    16'hfff9,
    16'hfff5,
    16'hfffc,
    16'hc,
    16'hfff1,
    16'hffff,
    16'h20,
    16'hfff4,
    16'hffdf,
    16'hffcc,
    16'hffd2,
    16'h6,
    16'hfff9,
    16'h35,
    16'h2,
    16'h17,
    16'hfffa,
    16'h0,
    16'h5,
    16'h2c,
    16'h23,
    16'h27,
    16'hc,
    16'h6,
    16'hfffa,
    16'hffeb,
    16'hffe2,
    16'hfff7,
    16'hfff5,
    16'he,
    16'hb,
    16'hffe7,
    16'hffe2,
    16'hffdd,
    16'hffed,
    16'hfffa,
    16'h13,
    16'h11,
    16'h42,
    16'h54,
    16'h21,
    16'h1c,
    16'hd,
    16'hfffc,
    16'h4,
    16'h10,
    16'h2f,
    16'h21,
    16'hffed,
    16'hfffb,
    16'hfff3,
    16'ha,
    16'h1c,
    16'h12,
    16'h4,
    16'h1c,
    16'hffdf,
    16'hc,
    16'h1b,
    16'h7,
    16'h1f,
    16'hffd1,
    16'hffee,
    16'hfffa,
    16'hffc5,
    16'hffe6,
    16'hfff5,
    16'hfff9,
    16'h47,
    16'h3c,
    16'hfffb,
    16'h14,
    16'h7,
    16'h1f,
    16'h7b,
    16'h35,
    16'h1b,
    16'h13,
    16'hfffe,
    16'hfff5,
    16'h1b,
    16'hffe4,
    16'hd,
    16'he,
    16'hfff5,
    16'h9,
    16'hfffd,
    16'hffff,
    16'h22,
    16'hfffe,
    16'h0,
    16'h13,
    16'hfff8,
    16'h5,
    16'hfff7,
    16'h16,
    16'he,
    16'h0,
    16'h3,
    16'hffef,
    16'ha,
    16'h0,
    16'hffd6,
    16'hffe5,
    16'hfffb,
    16'h14,
    16'hffdf,
    16'hfff0,
    16'h11,
    16'h8,
    16'hfffc,
    16'hfffe,
    16'h36,
    16'h2c,
    16'hffec,
    16'h28,
    16'hffe1,
    16'h9,
    16'he,
    16'h29,
    16'hfff3,
    16'h17,
    16'hffec,
    16'h1a,
    16'hfffd,
    16'hffe9,
    16'h3,
    16'h11,
    16'hffef,
    16'h15,
    16'hffe0,
    16'h3,
    16'hc,
    16'hffe4,
    16'h3,
    16'hffed,
    16'h13,
    16'h2,
    16'hffd9,
    16'hffbe,
    16'hfff9,
    16'hffe7,
    16'hffff,
    16'h8,
    16'h15,
    16'hf,
    16'hfff1,
    16'he,
    16'h3b,
    16'h40,
    16'hfffb,
    16'hb,
    16'h28,
    16'hfffd,
    16'h37,
    16'hfff2,
    16'hfffa,
    16'h18,
    16'hffff,
    16'h11,
    16'h3c,
    16'h16,
    16'hfff9,
    16'h0,
    16'hffe5,
    16'h4,
    16'hffef,
    16'h1,
    16'hffc8,
    16'hffd5,
    16'hffd2,
    16'hffdc,
    16'hffc5,
    16'hffe7,
    16'h11,
    16'hfff6,
    16'hffe2,
    16'hffcc,
    16'hffea,
    16'hfff0,
    16'h3,
    16'hfff5,
    16'h11,
    16'hffe8,
    16'hffe4,
    16'h14,
    16'h9,
    16'hffee,
    16'h8,
    16'hc,
    16'hffff,
    16'hffe4,
    16'h11,
    16'h10,
    16'h19,
    16'h21,
    16'hfffd,
    16'hfffd,
    16'hfff4,
    16'hffe3,
    16'hffdc,
    16'h9,
    16'h13,
    16'hfffe,
    16'hffe7,
    16'hfff5,
    16'hfff7,
    16'hc,
    16'he,
    16'hfff3,
    16'hffee,
    16'hffe6,
    16'hffef,
    16'hfffb,
    16'hffec,
    16'hfff4,
    16'h18,
    16'hffef,
    16'hffe2,
    16'hffbd,
    16'hfff6,
    16'h15,
    16'h2,
    16'h21,
    16'hfff9,
    16'hffeb,
    16'hffdb,
    16'hffde,
    16'h17,
    16'h11,
    16'hfff8,
    16'h9,
    16'hfffc,
    16'hd,
    16'h23,
    16'hfff5,
    16'ha,
    16'ha,
    16'hfff8,
    16'h6,
    16'hfff3,
    16'hfffb,
    16'hffed,
    16'hfff4,
    16'h7,
    16'hfff7,
    16'hffe3,
    16'hffe7,
    16'hffff,
    16'h13,
    16'hfff9,
    16'hf,
    16'h9,
    16'ha,
    16'h5,
    16'h31,
    16'h33,
    16'h1e,
    16'hfffd,
    16'h5,
    16'h0,
    16'hffc5,
    16'hffdf,
    16'hffe8,
    16'h14,
    16'hffd1,
    16'h1a,
    16'hffd9,
    16'h6,
    16'hfff9,
    16'hfff6,
    16'hfffb,
    16'h1f,
    16'hffec,
    16'hffee,
    16'h1,
    16'he,
    16'h33,
    16'h8,
    16'h15,
    16'h4,
    16'h10,
    16'hffe4,
    16'hfffc,
    16'hffe6,
    16'h5,
    16'hfffd,
    16'hffe8,
    16'h4,
    16'h10,
    16'h6,
    16'h15,
    16'hffe7,
    16'hf,
    16'hfff8,
    16'h1,
    16'h10,
    16'h14,
    16'hd,
    16'hfff4,
    16'h13,
    16'h8,
    16'h16,
    16'he,
    16'h6,
    16'h16,
    16'hffea,
    16'hffdf,
    16'hffe6,
    16'h0,
    16'hfffc,
    16'h7,
    16'h10,
    16'h14,
    16'hfff2,
    16'hffe8,
    16'hfff6,
    16'h3,
    16'h2,
    16'h8,
    16'hffef,
    16'hffd0,
    16'hffd2,
    16'hfff0,
    16'hfff4,
    16'hffef,
    16'hffd9,
    16'h3,
    16'hfffd,
    16'hfffa,
    16'h3,
    16'h6,
    16'hfff4,
    16'hffe5,
    16'h8,
    16'h1b,
    16'hffee,
    16'hffd8,
    16'hffeb,
    16'hfff1,
    16'h25,
    16'hffef,
    16'h11,
    16'h18,
    16'hfff8,
    16'h3,
    16'hd,
    16'h18,
    16'h1,
    16'h5,
    16'h17,
    16'h1b,
    16'h1a,
    16'h5,
    16'h3,
    16'h19,
    16'hfff8,
    16'h11,
    16'hb,
    16'hc,
    16'h4,
    16'h17,
    16'h27,
    16'h1f,
    16'h8,
    16'hffea,
    16'h2,
    16'hfff6,
    16'hfff6,
    16'hffda,
    16'hffd4,
    16'hffff,
    16'hfff5,
    16'hffdd,
    16'hffc2,
    16'hffd2,
    16'hffd7,
    16'h6,
    16'hfff4,
    16'h3,
    16'h27,
    16'hfffc,
    16'h13,
    16'h12,
    16'hfff6,
    16'hc,
    16'hd,
    16'h15,
    16'h1d,
    16'hc,
    16'h2,
    16'h10,
    16'h15,
    16'h2c,
    16'h4,
    16'hfff9,
    16'hffe4,
    16'hffe6,
    16'hffeb,
    16'ha,
    16'hf,
    16'h16,
    16'h16,
    16'h5,
    16'h18,
    16'hffe7,
    16'hfffd,
    16'h11,
    16'hfff8,
    16'hfffa,
    16'hffea,
    16'hffed,
    16'hffef,
    16'h16,
    16'hffe9,
    16'hfff6,
    16'ha,
    16'hffd9,
    16'h0,
    16'h9,
    16'hffe8,
    16'hfffa,
    16'h16,
    16'h18,
    16'hfff9,
    16'h8,
    16'h6,
    16'h2,
    16'hfffb,
    16'hffeb,
    16'h0,
    16'h12,
    16'h0,
    16'hfff6,
    16'h3,
    16'hd,
    16'h27,
    16'hc,
    16'hffef,
    16'h1d,
    16'h55,
    16'h33,
    16'h3b,
    16'h5,
    16'hfffd,
    16'h2d,
    16'h13,
    16'hfff1,
    16'h36,
    16'hffda,
    16'hfff9,
    16'h16,
    16'hffe5,
    16'h13,
    16'hf,
    16'hffee,
    16'h12,
    16'hc,
    16'hfff4,
    16'h23,
    16'h3,
    16'hfff5,
    16'h1,
    16'hfff3,
    16'hfff2,
    16'he,
    16'h2,
    16'hf,
    16'h15,
    16'h3,
    16'h0,
    16'h20,
    16'h6,
    16'hfffd,
    16'h9,
    16'hd,
    16'h32,
    16'h22,
    16'hfff3,
    16'hfffc,
    16'h13,
    16'h1,
    16'hffcb,
    16'hfffe,
    16'hffd3,
    16'hfff4,
    16'hfff5,
    16'hfffc,
    16'h5,
    16'hffe1,
    16'hffe9,
    16'hffff,
    16'hffee,
    16'h14,
    16'h1b,
    16'h1e,
    16'h1c,
    16'h5,
    16'hfff5,
    16'h19,
    16'h13,
    16'h17,
    16'h14,
    16'hd,
    16'hffed,
    16'h3,
    16'hffe8,
    16'h10,
    16'hfff7,
    16'h13,
    16'hfff3,
    16'h4,
    16'hff8f,
    16'hff8b,
    16'hffa7,
    16'h9,
    16'hfffd,
    16'hfffd,
    16'hff9a,
    16'hffc4,
    16'hffba,
    16'hfff4,
    16'ha,
    16'h2b,
    16'hf,
    16'h1f,
    16'h32,
    16'hfff9,
    16'hffec,
    16'hfff8,
    16'hd,
    16'h27,
    16'h27,
    16'hfff6,
    16'hffff,
    16'hffc2,
    16'hffab,
    16'hffd2,
    16'hffef,
    16'h4,
    16'h12,
    16'hfff0,
    16'h13,
    16'hfffd,
    16'h0,
    16'hfff0,
    16'h2,
    16'h3,
    16'h3,
    16'hfff8,
    16'h2,
    16'hfff9,
    16'h15,
    16'hf,
    16'hffff,
    16'hc,
    16'h24,
    16'h8,
    16'hfff5,
    16'h8,
    16'h11,
    16'h19,
    16'he,
    16'h19,
    16'hfff5,
    16'h12,
    16'h14,
    16'hfff6,
    16'hfff0,
    16'hfff4,
    16'hfffa,
    16'hfff0,
    16'h10,
    16'h10,
    16'h13,
    16'hffef,
    16'hfff4,
    16'h1,
    16'hfff4,
    16'h12,
    16'hfff0,
    16'hfff1,
    16'hfffb,
    16'h35,
    16'h1a,
    16'hffe1,
    16'hffb8,
    16'hffe1,
    16'hfff1,
    16'h35,
    16'h22,
    16'hffd8,
    16'hffcc,
    16'hffd9,
    16'hfff1,
    16'hfff6,
    16'hffef,
    16'hfffc,
    16'h1d,
    16'ha,
    16'hffe8,
    16'hffe8,
    16'hffee,
    16'hfffb,
    16'hf,
    16'h5,
    16'hffff,
    16'hffef,
    16'h13,
    16'hfffe,
    16'h10,
    16'hfff6,
    16'hfffe,
    16'h3,
    16'hfffe,
    16'hffff,
    16'h38,
    16'h2c,
    16'hfff4,
    16'hfff1,
    16'hffec,
    16'h1,
    16'h12,
    16'h45,
    16'hfff7,
    16'h0,
    16'hfffb,
    16'hffdd,
    16'hffa3,
    16'hfff5,
    16'hd,
    16'hffff,
    16'hfffa,
    16'hffdd,
    16'hffd5,
    16'hffe5,
    16'h12,
    16'h1,
    16'hfff7,
    16'h16,
    16'h8,
    16'h14,
    16'h12,
    16'h8,
    16'hffeb,
    16'h7,
    16'h1e,
    16'hfff1,
    16'h4,
    16'h2,
    16'hffea,
    16'hffee,
    16'hffe5,
    16'hfff8,
    16'hfff8,
    16'hffde,
    16'h9,
    16'h15,
    16'hf,
    16'h43,
    16'h8,
    16'h2,
    16'hfff1,
    16'hfffe,
    16'h15,
    16'h2a,
    16'h2,
    16'ha,
    16'hffed,
    16'h2e,
    16'hffdd,
    16'hffd0,
    16'h14,
    16'he,
    16'h8,
    16'h9,
    16'hffe3,
    16'hffdd,
    16'h14,
    16'h1c,
    16'hb,
    16'hfff2,
    16'h14,
    16'hfffe,
    16'hffee,
    16'hffee,
    16'hfff3,
    16'h9,
    16'h12,
    16'h40,
    16'hffe4,
    16'hffec,
    16'hfffe,
    16'h20,
    16'h1c,
    16'h36,
    16'hfff3,
    16'h1d,
    16'h2a,
    16'hfff4,
    16'h33,
    16'h54,
    16'h1c,
    16'hfffa,
    16'he,
    16'h19,
    16'hfffb,
    16'h1,
    16'h35,
    16'h1d,
    16'h6,
    16'hc,
    16'hffdd,
    16'hffe8,
    16'hf,
    16'h23,
    16'h0,
    16'h12,
    16'hffde,
    16'hffef,
    16'hfff6,
    16'hfffe,
    16'hfff9,
    16'hfff4,
    16'h28,
    16'h3,
    16'hfff1,
    16'hfff5,
    16'h22,
    16'hffe4,
    16'hffb2,
    16'hffdc,
    16'hfff9,
    16'hfff8,
    16'hfffe,
    16'he,
    16'hffdb,
    16'hffe5,
    16'h19,
    16'hffea,
    16'hfff3,
    16'hfff8,
    16'h12,
    16'h1,
    16'hffff,
    16'h28,
    16'h19,
    16'h12,
    16'ha,
    16'h7,
    16'h4,
    16'h7,
    16'h1d,
    16'h2c,
    16'h5,
    16'hffea,
    16'hffef,
    16'h5,
    16'hfff3,
    16'hfff4,
    16'h12,
    16'hfffc,
    16'hfffa,
    16'hffe9,
    16'h1a,
    16'h9,
    16'h1e,
    16'h1a,
    16'hffec,
    16'ha,
    16'hfffb,
    16'h12,
    16'h17,
    16'hfff5,
    16'h1a,
    16'hfff4,
    16'hfffa,
    16'hffe9,
    16'hffe9,
    16'hfff4,
    16'hfff5,
    16'hfff4,
    16'hfff1,
    16'hfffc,
    16'h3,
    16'hb,
    16'h9,
    16'h7,
    16'hd,
    16'hfff3,
    16'h19,
    16'hffeb,
    16'hfff4,
    16'hfff6,
    16'h0,
    16'hfff3,
    16'h1b,
    16'hfff5,
    16'hfffe,
    16'hfff9,
    16'h3,
    16'hfffb,
    16'hc,
    16'h2e,
    16'hffe8,
    16'hfffd,
    16'h20,
    16'h16,
    16'h20,
    16'h19,
    16'hfff9,
    16'hfffa,
    16'hf,
    16'h10,
    16'h3,
    16'hfffa,
    16'h13,
    16'hfff1,
    16'h1,
    16'hfff8,
    16'hfffa,
    16'h4,
    16'hffe4,
    16'h8,
    16'h1c,
    16'ha,
    16'hc,
    16'hf,
    16'h4,
    16'hfff9,
    16'h12,
    16'h8,
    16'h15,
    16'hfff7,
    16'hffd4,
    16'hffd5,
    16'hffed,
    16'h4,
    16'hfff6,
    16'h2c,
    16'hffe0,
    16'hffd8,
    16'hffea,
    16'h10,
    16'h1a,
    16'h7,
    16'h17,
    16'h27,
    16'hfffe,
    16'h16,
    16'hfffb,
    16'hffe5,
    16'hfff4,
    16'h30,
    16'h33,
    16'hfffa,
    16'hffe2,
    16'h3,
    16'he,
    16'hf,
    16'h27,
    16'h11,
    16'h14,
    16'ha,
    16'h15,
    16'he,
    16'hfff7,
    16'h11,
    16'hfff2,
    16'hfff6,
    16'hb,
    16'hfff4,
    16'hfffb,
    16'hffef,
    16'hffe7,
    16'hffe9,
    16'hfff0,
    16'hffd3,
    16'hffe9,
    16'hffcf,
    16'he,
    16'hffd1,
    16'hffef,
    16'hffec,
    16'hfffe,
    16'h1,
    16'hfffb,
    16'h7,
    16'h13,
    16'h9,
    16'h14,
    16'hb,
    16'hb,
    16'h1a,
    16'h1f,
    16'h16,
    16'h18,
    16'hffff,
    16'ha,
    16'h8,
    16'h8,
    16'hffee,
    16'hfff0,
    16'h14,
    16'h13,
    16'hfffe,
    16'hffe3,
    16'he,
    16'hffef,
    16'hfff0,
    16'h15,
    16'h5,
    16'hfff9,
    16'h5,
    16'h0,
    16'hfff9,
    16'hffd5,
    16'hffdd,
    16'hfffe,
    16'hfffa,
    16'h11,
    16'he,
    16'hfffe,
    16'hfff1,
    16'h4,
    16'hfffe,
    16'hffd5,
    16'hffeb,
    16'hd,
    16'hfffe,
    16'h1,
    16'ha,
    16'hfffb,
    16'h1,
    16'hfff3,
    16'hfff6,
    16'hfff5,
    16'hffee,
    16'h1,
    16'ha,
    16'h12,
    16'hfffd,
    16'hfff1,
    16'hfff0,
    16'hffff,
    16'h36,
    16'h5a,
    16'h16,
    16'h11,
    16'hffff,
    16'hfffc,
    16'h4f,
    16'h53,
    16'h26,
    16'h7,
    16'h3e,
    16'h2d,
    16'h1d,
    16'h9,
    16'hfff3,
    16'hfff5,
    16'h28,
    16'h11,
    16'hfffe,
    16'hfffa,
    16'hffed,
    16'hffff,
    16'h1f,
    16'hfffc,
    16'hfff5,
    16'hc,
    16'hfffd,
    16'hfffc,
    16'hb,
    16'h10,
    16'hfffc,
    16'hffec,
    16'h2,
    16'h2,
    16'h7,
    16'hfff2,
    16'h13,
    16'h3c,
    16'h9,
    16'h12,
    16'h5,
    16'h8,
    16'h2b,
    16'h22,
    16'hd,
    16'h8,
    16'h9,
    16'h2f,
    16'h1e,
    16'hfff3,
    16'hffec,
    16'h1a,
    16'h10,
    16'hfffa,
    16'h7,
    16'h10,
    16'hffea,
    16'hffeb,
    16'hc,
    16'ha,
    16'hffec,
    16'h18,
    16'he,
    16'hffed,
    16'hfff8,
    16'h2,
    16'hffdc,
    16'hffd4,
    16'hfff1,
    16'h17,
    16'h7,
    16'h1f,
    16'hffd0,
    16'hff99,
    16'hffb0,
    16'hd,
    16'h14,
    16'hf,
    16'hffea,
    16'hffd9,
    16'hffaf,
    16'hffec,
    16'hffe1,
    16'hffdc,
    16'hffde,
    16'h25,
    16'h1c,
    16'hfffb,
    16'hffee,
    16'hffef,
    16'hfffc,
    16'h29,
    16'h15,
    16'h10,
    16'h5,
    16'hffe8,
    16'hffea,
    16'hfffe,
    16'h1d,
    16'h6,
    16'h10,
    16'hffe9,
    16'hffef,
    16'hfff4,
    16'hb,
    16'hfffc,
    16'hffe7,
    16'hffeb,
    16'h14,
    16'h1a,
    16'h15,
    16'hfff1,
    16'h9,
    16'hffee,
    16'h2e,
    16'h40,
    16'h50,
    16'hfff9,
    16'h23,
    16'h1e,
    16'h38,
    16'h6,
    16'h2,
    16'h19,
    16'h14,
    16'hf,
    16'h7,
    16'hffff,
    16'hffea,
    16'h4,
    16'h12,
    16'hfff5,
    16'hffea,
    16'hfff0,
    16'h15,
    16'hffeb,
    16'hffe6,
    16'hffe7,
    16'hfff5,
    16'h9,
    16'hffe6,
    16'hffec,
    16'h13,
    16'hfffa,
    16'h1e,
    16'h27,
    16'h32,
    16'hb,
    16'h22,
    16'h6,
    16'h33,
    16'h59,
    16'h8a,
    16'h3,
    16'h2b,
    16'h36,
    16'h27,
    16'h7,
    16'hffe3,
    16'h1,
    16'h0,
    16'hd,
    16'hfffe,
    16'hfff8,
    16'h6,
    16'hffff,
    16'hf,
    16'h9,
    16'hd,
    16'hfff1,
    16'hfff5,
    16'h14,
    16'h3,
    16'hfff2,
    16'hffed,
    16'hffe9,
    16'hfffc,
    16'hfff8,
    16'h10,
    16'hfffc,
    16'hffea,
    16'hfff1,
    16'hffef,
    16'h3,
    16'hb,
    16'hfff1,
    16'hfff7,
    16'hd,
    16'he,
    16'hfff7,
    16'hffe2,
    16'hfff6,
    16'hfffe,
    16'h1,
    16'hffe3,
    16'hfff1,
    16'h11,
    16'hfff8,
    16'h8,
    16'h2,
    16'hfff9,
    16'hfff0,
    16'h8,
    16'hffe8,
    16'hfff1,
    16'hfff6,
    16'h16,
    16'hf,
    16'h17,
    16'hfffb,
    16'hfff8,
    16'hfff8,
    16'h10,
    16'h15,
    16'hfff9,
    16'hffd3,
    16'hffc6,
    16'hffbc,
    16'h2,
    16'hffef,
    16'h19,
    16'h1,
    16'hffcb,
    16'hfff2,
    16'h19,
    16'hffe1,
    16'h2d,
    16'h1f,
    16'h4,
    16'h27,
    16'hc,
    16'hfff7,
    16'h21,
    16'h2e,
    16'h25,
    16'hc,
    16'hffe5,
    16'hffeb,
    16'hffef,
    16'hffe3,
    16'hfff5,
    16'h4,
    16'h2,
    16'h17,
    16'h14,
    16'h18,
    16'h18,
    16'h32,
    16'h20,
    16'hfffb,
    16'hffde,
    16'hfff6,
    16'h11,
    16'h8,
    16'hffe5,
    16'hfff6,
    16'hfff7,
    16'h7,
    16'hfff8,
    16'hfff5,
    16'hffff,
    16'h5,
    16'hffff,
    16'he,
    16'ha,
    16'h6,
    16'h3,
    16'hffff,
    16'h13,
    16'h15,
    16'h8,
    16'h22,
    16'h14,
    16'hffee,
    16'h2c,
    16'hfffb,
    16'hffb3,
    16'hffde,
    16'hf,
    16'h14,
    16'h9,
    16'hfff2,
    16'hffff,
    16'hffe4,
    16'hffe7,
    16'hffdd,
    16'hfff0,
    16'h8,
    16'hffe2,
    16'h22,
    16'h45,
    16'hffdd,
    16'hffe4,
    16'hffef,
    16'hfffc,
    16'h1f,
    16'hfffe,
    16'hffe8,
    16'hffd9,
    16'hfff4,
    16'h19,
    16'hfff6,
    16'hffdc,
    16'hfff6,
    16'h0,
    16'hfffa,
    16'h10,
    16'h19,
    16'h12,
    16'hfff6,
    16'ha,
    16'h27,
    16'hfff3,
    16'h11,
    16'h7,
    16'hc,
    16'hffe8,
    16'h4,
    16'hfff8,
    16'hfff7,
    16'hffec,
    16'hfff9,
    16'hffd9,
    16'hfff0,
    16'hffe9,
    16'h17,
    16'hf,
    16'hffda,
    16'h19,
    16'h19,
    16'h2,
    16'hf,
    16'h12,
    16'hffec,
    16'hffe9,
    16'hd,
    16'ha,
    16'hf,
    16'hfffc,
    16'h0,
    16'h1d,
    16'hfff2,
    16'hc,
    16'hfff3,
    16'hffef,
    16'hfff4,
    16'h8,
    16'h3,
    16'h2a,
    16'h16,
    16'h7,
    16'h3,
    16'hfff7,
    16'hfff3,
    16'h0,
    16'hffe5,
    16'hffee,
    16'hffd9,
    16'hfffc,
    16'h22,
    16'h7,
    16'hffaf,
    16'hffe1,
    16'hfff7,
    16'h0,
    16'hfff9,
    16'h9,
    16'hffe8,
    16'h11,
    16'hffe8,
    16'hf,
    16'h15,
    16'h4,
    16'h12,
    16'hfff4,
    16'hffcd,
    16'hfffd,
    16'h1c,
    16'h2e,
    16'h20,
    16'h1,
    16'h11,
    16'hfff9,
    16'hffe4,
    16'hffe7,
    16'hffdd,
    16'h3,
    16'h13,
    16'hffef,
    16'h17,
    16'hffe7,
    16'hffe8,
    16'hb,
    16'h6,
    16'hffe8,
    16'h28,
    16'h2,
    16'he,
    16'hffeb,
    16'hffe9,
    16'hffec,
    16'hc,
    16'h27,
    16'hffee,
    16'hffef,
    16'hfff1,
    16'hffee,
    16'hfff3,
    16'hffdc,
    16'h0,
    16'h6,
    16'hffe6,
    16'hfffb,
    16'hfff3,
    16'hfffe,
    16'hb,
    16'h15,
    16'hfff8,
    16'hffe5,
    16'h11,
    16'h7,
    16'hfff5,
    16'h10,
    16'h2,
    16'h0,
    16'hfff7,
    16'hffe5,
    16'hffe1,
    16'hfff7,
    16'h8,
    16'h7,
    16'hffed,
    16'hffc4,
    16'hffea,
    16'hfffa,
    16'h5,
    16'h3,
    16'hffe8,
    16'hfffd,
    16'h1d,
    16'h3a,
    16'hf,
    16'hf,
    16'h7,
    16'hc,
    16'h1e,
    16'hfff8,
    16'hfffc,
    16'h1a,
    16'hfff5,
    16'h25,
    16'hffff,
    16'h1,
    16'hffdb,
    16'hffcc,
    16'hffcc,
    16'hffd2,
    16'hfff5,
    16'hfffd,
    16'hfffc,
    16'hfff9,
    16'h19,
    16'h10,
    16'h2,
    16'hb,
    16'h11,
    16'ha,
    16'h1,
    16'ha,
    16'h4,
    16'h12,
    16'hffec,
    16'hfff3,
    16'hfffa,
    16'h0,
    16'hfff9,
    16'hc,
    16'hffd3,
    16'hffb5,
    16'h0,
    16'hfff1,
    16'ha,
    16'hfff2,
    16'hfff8,
    16'hffc2,
    16'hffed,
    16'hfff3,
    16'hfffc,
    16'h23,
    16'h11,
    16'hfff1,
    16'h2b,
    16'hb,
    16'ha,
    16'hffed,
    16'hfff4,
    16'hfffc,
    16'hffe7,
    16'h17,
    16'hffe8,
    16'hfff0,
    16'hffea,
    16'ha,
    16'h2e,
    16'h11,
    16'hffe6,
    16'hffee,
    16'h4,
    16'hd,
    16'h32,
    16'h2e,
    16'hfff1,
    16'hfff3,
    16'hffc9,
    16'hffd8,
    16'h3,
    16'hfff5,
    16'hd,
    16'hfffc,
    16'ha,
    16'hffb9,
    16'hffd0,
    16'hffe6,
    16'hffef,
    16'h0,
    16'h1f,
    16'h14,
    16'h20,
    16'h3f,
    16'h4,
    16'h18,
    16'h2,
    16'h1a,
    16'h31,
    16'h43,
    16'h4e,
    16'h1f,
    16'hfff8,
    16'hffff,
    16'hfffb,
    16'h1c,
    16'hfffb,
    16'hffe8,
    16'hfff5,
    16'h1,
    16'hffec,
    16'hffed,
    16'hffca,
    16'hfff8,
    16'h15,
    16'h14,
    16'hffeb,
    16'hd,
    16'hfff8,
    16'hb,
    16'hc,
    16'h10,
    16'h18,
    16'h1c,
    16'h1a,
    16'h20,
    16'h6,
    16'hffe8,
    16'hfff1,
    16'hffeb,
    16'h18,
    16'h0,
    16'h12,
    16'hffef,
    16'hffed,
    16'hffd8,
    16'hffdb,
    16'hfff1,
    16'h1,
    16'hffee,
    16'hffe3,
    16'hfff7,
    16'h41,
    16'h36,
    16'he,
    16'hffdd,
    16'hffc3,
    16'hfff5,
    16'h1d,
    16'hffe5,
    16'hfff4,
    16'hffc0,
    16'hffcd,
    16'hffe3,
    16'hfff2,
    16'hffe4,
    16'h1c,
    16'hfffd,
    16'hffff,
    16'hffe7,
    16'hfff4,
    16'h15,
    16'hb,
    16'ha,
    16'hfffe,
    16'h1b,
    16'hfff7,
    16'hf,
    16'hffe5,
    16'hffea,
    16'h11,
    16'h3,
    16'hffef,
    16'hfff7,
    16'hfffc,
    16'hfffb,
    16'h0,
    16'h17,
    16'h13,
    16'h1d,
    16'h4,
    16'h2,
    16'hffe3,
    16'h8,
    16'hfff3,
    16'hffe3,
    16'hffe9,
    16'h5,
    16'hffd2,
    16'hffd4,
    16'hffec,
    16'hffec,
    16'h0,
    16'h3,
    16'hffe9,
    16'h6,
    16'h10,
    16'hffeb,
    16'hffe6,
    16'hffec,
    16'hffef,
    16'hfffd,
    16'hfff9,
    16'h12,
    16'hfffc,
    16'hfffc,
    16'h34,
    16'h28,
    16'h12,
    16'h23,
    16'h9,
    16'h11,
    16'h3d,
    16'hfff2,
    16'hffb0,
    16'hffe3,
    16'h17,
    16'h1e,
    16'h1b,
    16'hffec,
    16'hffb4,
    16'h22,
    16'hfff1,
    16'h16,
    16'h28,
    16'h0,
    16'h17,
    16'h38,
    16'hc,
    16'hfff5,
    16'hc,
    16'hffde,
    16'h9,
    16'hfff5,
    16'hffe9,
    16'ha,
    16'hffea,
    16'hfff4,
    16'hfffd,
    16'hffe2,
    16'h9,
    16'h7,
    16'h0,
    16'hfffc,
    16'hffc5,
    16'hffe2,
    16'h16,
    16'h8,
    16'h20,
    16'h1d,
    16'h38,
    16'h23,
    16'hffed,
    16'hffea,
    16'hfff0,
    16'hffff,
    16'h10,
    16'h4,
    16'h14,
    16'hffd2,
    16'hffd5,
    16'hffed,
    16'hffe1,
    16'hffe8,
    16'hffec,
    16'hffe9,
    16'hffcf,
    16'hffdd,
    16'h3,
    16'hfffe,
    16'hc,
    16'hfffb,
    16'h19,
    16'hfff5,
    16'hc,
    16'h16,
    16'hb,
    16'ha,
    16'h22,
    16'h7,
    16'hffff,
    16'h6,
    16'hffef,
    16'hffef,
    16'hffaf,
    16'hffc8,
    16'h1b,
    16'h22,
    16'hfff6,
    16'hffed,
    16'hffbc,
    16'hffcd,
    16'h12,
    16'hffdc,
    16'h8,
    16'h6,
    16'hffec,
    16'hfff5,
    16'h1c,
    16'hd,
    16'h7,
    16'h2a,
    16'hfffa,
    16'h0,
    16'he,
    16'h13,
    16'hffe0,
    16'hffff,
    16'h39,
    16'h25,
    16'hd,
    16'hfff0,
    16'h7,
    16'hd,
    16'hffee,
    16'hfffd,
    16'h18,
    16'hfffe,
    16'he,
    16'h1f,
    16'h25,
    16'h7,
    16'h2,
    16'he,
    16'hfff5,
    16'h1b,
    16'h10,
    16'hfffb,
    16'h13,
    16'hfff4,
    16'h1b,
    16'h3,
    16'hfff7,
    16'hffe9,
    16'hf,
    16'hfffc,
    16'h5,
    16'hfffa,
    16'hffeb,
    16'h6,
    16'he,
    16'he,
    16'h11,
    16'hfff3,
    16'hfffd,
    16'hfffe,
    16'hfff4,
    16'hffec,
    16'h9,
    16'hfff6,
    16'hffe1,
    16'h6,
    16'h7,
    16'h13,
    16'hffee,
    16'h27,
    16'h19,
    16'h1f,
    16'hfffc,
    16'hffe8,
    16'hb,
    16'h4,
    16'hffc6,
    16'h2f,
    16'h22,
    16'h4,
    16'h5,
    16'hffcf,
    16'hffc5,
    16'hfffd,
    16'h4,
    16'hffea,
    16'hfff1,
    16'hffe6,
    16'hffea,
    16'hffe7,
    16'hffe7,
    16'hffea,
    16'hfff3,
    16'hfffa,
    16'hf,
    16'h23,
    16'h0,
    16'h2,
    16'h4,
    16'hfffd,
    16'hffe5,
    16'hffdf,
    16'hffe7,
    16'h3,
    16'h11,
    16'h16,
    16'hfff5,
    16'hfffa,
    16'h2f,
    16'h33,
    16'hfffb,
    16'hfff9,
    16'h9,
    16'hffdb,
    16'hfffa,
    16'hb,
    16'h9,
    16'hffeb,
    16'hffdc,
    16'h31,
    16'h1c,
    16'h4,
    16'h7,
    16'hfff7,
    16'hfff0,
    16'h1f,
    16'hffdb,
    16'hffee,
    16'hffc3,
    16'hffe4,
    16'h3b,
    16'hfff6,
    16'hffd4,
    16'he,
    16'h15,
    16'h4,
    16'hfffb,
    16'hffd9,
    16'hfff4,
    16'h6,
    16'h3d,
    16'h2b,
    16'ha,
    16'hfffb,
    16'h1d,
    16'hffe4,
    16'h20,
    16'h1f,
    16'hffec,
    16'h14,
    16'hfff3,
    16'h21,
    16'h12,
    16'hfff5,
    16'hfffb,
    16'h8,
    16'h17,
    16'h18,
    16'h4,
    16'h3,
    16'hffe1,
    16'hd,
    16'h1b,
    16'hfffe,
    16'hffd4,
    16'hffd3,
    16'hfffd,
    16'h16,
    16'hffb2,
    16'hffcb,
    16'h1a,
    16'h17,
    16'hffeb,
    16'hfff2,
    16'hd,
    16'hfff6,
    16'h14,
    16'h24,
    16'h23,
    16'hfffc,
    16'hfff3,
    16'hffd1,
    16'h1b,
    16'h9,
    16'h0,
    16'hc,
    16'hffef,
    16'hffe1,
    16'h16,
    16'hffed,
    16'hffc9,
    16'h1b,
    16'hffe2,
    16'hffea,
    16'h4,
    16'hffff,
    16'hffe4,
    16'hffd7,
    16'h5,
    16'h4,
    16'h3,
    16'hffd6,
    16'hfff4,
    16'hffb2,
    16'hffde,
    16'h0,
    16'h19,
    16'ha,
    16'hfff6,
    16'hffed,
    16'hfff0,
    16'hffe8,
    16'h18,
    16'h24,
    16'h9,
    16'h19,
    16'h1d,
    16'hfff3,
    16'hfff8,
    16'hfffa,
    16'hffdc,
    16'hfff0,
    16'hb,
    16'h15,
    16'hffe9,
    16'hffe6,
    16'hffcc,
    16'h1b,
    16'h5,
    16'hfffc,
    16'ha,
    16'hffe2,
    16'hfff9,
    16'hfff0,
    16'hffca,
    16'hffd9,
    16'h18,
    16'h48,
    16'h34,
    16'h17,
    16'hfff1,
    16'hffe2,
    16'hfffe,
    16'h7,
    16'hf,
    16'hf,
    16'hfff9,
    16'hfff5,
    16'hfffc,
    16'hfff5,
    16'h10,
    16'h14,
    16'h0,
    16'h0,
    16'hfffc,
    16'hfff5,
    16'hfff9,
    16'hffdd,
    16'hfffa,
    16'hb,
    16'hfffc,
    16'h22,
    16'h13,
    16'h11,
    16'hffee,
    16'hffea,
    16'h3,
    16'hfff4,
    16'h3,
    16'h4,
    16'h12,
    16'hffee,
    16'h1,
    16'hc,
    16'hfffa,
    16'h2,
    16'hfff2,
    16'h1a,
    16'hffea,
    16'h12,
    16'h10,
    16'hffeb,
    16'ha,
    16'hfffb,
    16'h1d,
    16'h28,
    16'h17,
    16'hf,
    16'h15,
    16'ha,
    16'h1,
    16'h0,
    16'hffe2,
    16'h2,
    16'h7,
    16'h1,
    16'h4,
    16'hffff,
    16'hffee,
    16'hffe5,
    16'hfffe,
    16'h1,
    16'hffe6,
    16'he,
    16'hfffd,
    16'hffed,
    16'hffe4,
    16'hffed,
    16'h10,
    16'hffff,
    16'h1c,
    16'h20,
    16'hfffe,
    16'hffed,
    16'he,
    16'h4,
    16'h4,
    16'hfff3,
    16'hffe8,
    16'h13,
    16'hfff1,
    16'hfff0,
    16'h10,
    16'hffef,
    16'h18,
    16'hfff7,
    16'h2b,
    16'h25,
    16'h21,
    16'h18,
    16'h1e,
    16'hfff0,
    16'hfffc,
    16'h32,
    16'hffd8,
    16'hffc9,
    16'he,
    16'h15,
    16'h23,
    16'h14,
    16'hfff7,
    16'hffde,
    16'hfffd,
    16'h0,
    16'hfff0,
    16'hffe7,
    16'hffc7,
    16'hfff6,
    16'hfffe,
    16'hffe3,
    16'hffff,
    16'hffea,
    16'hfff8,
    16'hfff5,
    16'hfff2,
    16'hffee,
    16'hfff0,
    16'hfff2,
    16'hffd6,
    16'hc,
    16'h1c,
    16'h1f,
    16'h9,
    16'h18,
    16'hffd8,
    16'hffd8,
    16'h0,
    16'h8,
    16'hfff8,
    16'h1e,
    16'h44,
    16'hc,
    16'h2,
    16'hfff2,
    16'ha,
    16'h22,
    16'hfffb,
    16'hfff5,
    16'hfff4,
    16'he,
    16'h17,
    16'h25,
    16'h13,
    16'hfff9,
    16'h1a,
    16'hb,
    16'h0,
    16'h5,
    16'hffed,
    16'h1f,
    16'h10,
    16'hc,
    16'hfffb,
    16'h28,
    16'hfffa,
    16'hfff5,
    16'h15,
    16'hc,
    16'hfff5,
    16'h14,
    16'h14,
    16'h11,
    16'hfffc,
    16'h8,
    16'ha,
    16'hc,
    16'hd,
    16'h9,
    16'h1,
    16'hfffa,
    16'hfff2,
    16'h5,
    16'h20,
    16'h17,
    16'hb,
    16'h16,
    16'h15,
    16'hfff2,
    16'h19,
    16'h2b,
    16'hfff1,
    16'hffec,
    16'ha,
    16'hfff8,
    16'h1e,
    16'ha,
    16'h1d,
    16'hffff,
    16'h1,
    16'h1c,
    16'h2e,
    16'hffee,
    16'hffdd,
    16'h2,
    16'h8,
    16'h1c,
    16'h34,
    16'h1b,
    16'hfff7,
    16'hd,
    16'h18,
    16'h1c,
    16'hfffd,
    16'hffe9,
    16'h1b,
    16'h6,
    16'hfffc,
    16'hfffe,
    16'hfff2,
    16'h14,
    16'h16,
    16'h4,
    16'hffe8,
    16'hffef,
    16'hffe3,
    16'hfff0,
    16'ha,
    16'hfff4,
    16'h1a,
    16'hfff7,
    16'hfff8,
    16'hfff5,
    16'h15,
    16'hffea,
    16'hffff,
    16'h12,
    16'h14,
    16'h3,
    16'hffdf,
    16'hfff8,
    16'hfffa,
    16'hd,
    16'hfff7,
    16'h22,
    16'hffec,
    16'hfff7,
    16'h7,
    16'hfffd,
    16'h31,
    16'h20,
    16'hffff,
    16'h3,
    16'hffec,
    16'h19,
    16'hfff2,
    16'hfff5,
    16'h7,
    16'hfff6,
    16'h4,
    16'h14,
    16'h1,
    16'hf,
    16'h13,
    16'hfff9,
    16'h15,
    16'hffe1,
    16'hfff4,
    16'hffe0,
    16'hfff2,
    16'h4,
    16'h9,
    16'hffe7,
    16'hffeb,
    16'h3,
    16'h32,
    16'h9,
    16'hf,
    16'hb,
    16'h11,
    16'hfff3,
    16'h3b,
    16'ha,
    16'h11,
    16'h15,
    16'h24,
    16'hfffb,
    16'h18,
    16'hfff7,
    16'hfff6,
    16'h10,
    16'h9,
    16'h25,
    16'hffe9,
    16'hffd9,
    16'hd,
    16'hffee,
    16'h21,
    16'h3e,
    16'hc,
    16'hfff4,
    16'hfff3,
    16'h1b,
    16'h1,
    16'h8,
    16'h17,
    16'hfffe,
    16'hffe9,
    16'h7,
    16'hffef,
    16'hffe9,
    16'hffeb,
    16'hfff5,
    16'hc,
    16'h1d,
    16'h22,
    16'h5,
    16'hffec,
    16'h5,
    16'hfffd,
    16'hf,
    16'h2c,
    16'h21,
    16'hffe1,
    16'hfff7,
    16'h1f,
    16'h1d,
    16'h3,
    16'h20,
    16'h2a,
    16'h18,
    16'h6,
    16'hfff1,
    16'hffe1,
    16'hfff8,
    16'hfffd,
    16'hfff6,
    16'hffe5,
    16'hffe6,
    16'hfff6,
    16'hf,
    16'hb,
    16'h16,
    16'hf,
    16'hf,
    16'h1d,
    16'h12,
    16'hffe6,
    16'hffdd,
    16'h12,
    16'h15,
    16'h3a,
    16'h6b,
    16'h1d,
    16'hffff,
    16'hfff9,
    16'hfff9,
    16'hffcf,
    16'hffd1,
    16'h20,
    16'hffef,
    16'hffed,
    16'hffc5,
    16'hffba,
    16'hfff0,
    16'h1e,
    16'hfffe,
    16'hffe4,
    16'hffd1,
    16'hffd6,
    16'hffc8,
    16'hffb8,
    16'hffdf,
    16'h0,
    16'h11,
    16'hffe9,
    16'hfff0,
    16'h5,
    16'hffe9,
    16'h19,
    16'hd,
    16'hfff1,
    16'hfff2,
    16'hffe4,
    16'h8,
    16'hfff4,
    16'h4,
    16'hfffc,
    16'hfffa,
    16'hffe4,
    16'hffe3,
    16'hffee,
    16'hffea,
    16'hfffc,
    16'hfffc,
    16'he,
    16'hffe8,
    16'hffe9,
    16'hfffa,
    16'hfff1,
    16'hfff7,
    16'hfff5,
    16'hd,
    16'h8,
    16'hfff5,
    16'hb,
    16'hfffa,
    16'h1,
    16'h12,
    16'hffeb,
    16'hfff9,
    16'hfff1,
    16'hffed,
    16'hfffe,
    16'hfffa,
    16'h8,
    16'hfff4,
    16'hb,
    16'ha,
    16'h18,
    16'h1b,
    16'hffed,
    16'h27,
    16'h47,
    16'hb,
    16'hffe4,
    16'ha,
    16'hffe2,
    16'h2,
    16'h3b,
    16'he,
    16'h0,
    16'h2,
    16'hffea,
    16'h3,
    16'hf,
    16'h1,
    16'h12,
    16'h16,
    16'hd,
    16'h11,
    16'ha,
    16'hffff,
    16'hfffd,
    16'h8,
    16'hfffa,
    16'h2,
    16'hb,
    16'hc,
    16'h1,
    16'h10,
    16'hfffc,
    16'hffff,
    16'h5,
    16'hfffe,
    16'hfffb,
    16'h12,
    16'h8,
    16'h16,
    16'hffe2,
    16'hffee,
    16'h1c,
    16'h25,
    16'h5,
    16'hffe4,
    16'h1e,
    16'h8,
    16'hfff7,
    16'hffd5,
    16'hffee,
    16'h0,
    16'hffff,
    16'hffdd,
    16'hffdf,
    16'h3,
    16'h1d,
    16'h15,
    16'h11,
    16'h32,
    16'h35,
    16'he,
    16'h7,
    16'h9,
    16'hb,
    16'hb,
    16'h20,
    16'hb,
    16'h0,
    16'hffec,
    16'h5,
    16'hfff9,
    16'hd,
    16'h4,
    16'h6,
    16'hffda,
    16'hfff8,
    16'h7,
    16'h1d,
    16'h1a,
    16'hfff8,
    16'hffea,
    16'h3,
    16'h7,
    16'h1f,
    16'h22,
    16'hffe9,
    16'hffe8,
    16'h1,
    16'hfffe,
    16'hffd2,
    16'hffbb,
    16'hfffb,
    16'hfffc,
    16'hd,
    16'h1,
    16'h8,
    16'hd,
    16'h0,
    16'h1,
    16'h24,
    16'h13,
    16'hfffe,
    16'h7,
    16'hb,
    16'h1,
    16'h4,
    16'h1e,
    16'h28,
    16'h30,
    16'hffec,
    16'h10,
    16'hfffb,
    16'h10,
    16'hb,
    16'h8,
    16'h11,
    16'h16,
    16'hf,
    16'h7,
    16'h21,
    16'h11,
    16'hfff5,
    16'hfffa,
    16'hffea,
    16'h1c,
    16'h1a,
    16'hffff,
    16'hfff6,
    16'hfffa,
    16'h2e,
    16'h12,
    16'hfff2,
    16'hfffd,
    16'hffea,
    16'he,
    16'h12,
    16'h13,
    16'h21,
    16'hfffe,
    16'h22,
    16'hb,
    16'h21,
    16'h4,
    16'h13,
    16'h1e,
    16'hb,
    16'h7,
    16'h2c,
    16'h2e,
    16'h2,
    16'h0,
    16'hfffd,
    16'h17,
    16'h31,
    16'hfff5,
    16'h9,
    16'hfff9,
    16'hffe7,
    16'hffeb,
    16'h15,
    16'hd,
    16'h11,
    16'h2,
    16'h2,
    16'hfff9,
    16'h5,
    16'h18,
    16'h26,
    16'hfffb,
    16'hffee,
    16'hc,
    16'hffef,
    16'hffec,
    16'hffec,
    16'h0,
    16'h11,
    16'h2,
    16'hfffe,
    16'hfffb,
    16'hfffb,
    16'hffe8,
    16'hffe6,
    16'hfffb,
    16'hffd8,
    16'h34,
    16'hb,
    16'h11,
    16'hf,
    16'hffeb,
    16'hffd2,
    16'hffe6,
    16'h1,
    16'ha,
    16'hffec,
    16'h18,
    16'h14,
    16'hffe9,
    16'hffe1,
    16'h7,
    16'hffe7,
    16'hffeb,
    16'h14,
    16'hfff5,
    16'hffeb,
    16'hffed,
    16'hfffc,
    16'hfff8,
    16'h10,
    16'h28,
    16'h14,
    16'hfffe,
    16'h5,
    16'hfffa,
    16'hb,
    16'h1,
    16'hb,
    16'h18,
    16'h2,
    16'hffff,
    16'h1c,
    16'h17,
    16'hfff0,
    16'he,
    16'h9,
    16'hffe6,
    16'hfffb,
    16'hb,
    16'hc,
    16'he,
    16'he,
    16'h1,
    16'hffef,
    16'h1d,
    16'hfffe,
    16'hfff0,
    16'hfff8,
    16'hffe0,
    16'hffff,
    16'hffef,
    16'h2,
    16'hfff8,
    16'h17,
    16'hc,
    16'hfff6,
    16'hffff,
    16'h13,
    16'h3,
    16'h11,
    16'hffeb,
    16'hfff3,
    16'h22,
    16'h1d,
    16'h29,
    16'hfffc,
    16'hffef,
    16'hffe6,
    16'hffff,
    16'hfffc,
    16'h3,
    16'hc,
    16'h21,
    16'h24,
    16'h5,
    16'h19,
    16'h5,
    16'hffe4,
    16'hffbe,
    16'h4,
    16'hffff,
    16'hfff4,
    16'hffe0,
    16'hffee,
    16'hfff3,
    16'hfff7,
    16'hfffe,
    16'h4,
    16'h4,
    16'h16,
    16'hffef,
    16'he,
    16'h6,
    16'hfff9,
    16'hffeb,
    16'h17,
    16'hfff5,
    16'hffe6,
    16'hfffa,
    16'h10,
    16'h13,
    16'hfff9,
    16'hffc5,
    16'hffd2,
    16'h18,
    16'h3,
    16'ha,
    16'h13,
    16'hffff,
    16'h0,
    16'hffee,
    16'hfff7,
    16'h9,
    16'hfff8,
    16'hffef,
    16'hffd6,
    16'h10,
    16'h11,
    16'hffff,
    16'hfff3,
    16'hffcc,
    16'hffbc,
    16'hffd6,
    16'hffea,
    16'h14,
    16'hfffc,
    16'h5,
    16'hffea,
    16'hffe3,
    16'hffe4,
    16'hfff0,
    16'hffec,
    16'hfffc,
    16'h1d,
    16'h26,
    16'hb,
    16'hfffd,
    16'h11,
    16'hd,
    16'hffff,
    16'hfffc,
    16'hf,
    16'h25,
    16'hb,
    16'hffda,
    16'h9,
    16'h2d,
    16'h10,
    16'hfff8,
    16'ha,
    16'h2b,
    16'h54,
    16'h11,
    16'h0,
    16'hfffb,
    16'h1,
    16'hfff7,
    16'hd,
    16'hc,
    16'ha,
    16'hfff2,
    16'h15,
    16'h9,
    16'hfff0,
    16'hffed,
    16'hfffd,
    16'hfff3,
    16'hfff8,
    16'hffdd,
    16'hffe4,
    16'hffff,
    16'hffe8,
    16'hfff9,
    16'hc,
    16'h2,
    16'hffd3,
    16'hffc7,
    16'h2,
    16'hfff6,
    16'h10,
    16'hffdf,
    16'hffbf,
    16'hfffe,
    16'h10,
    16'hfffc,
    16'hfff0,
    16'hffc4,
    16'hffd6,
    16'hffe0,
    16'hffe0,
    16'hfffd,
    16'h6,
    16'h23,
    16'h15,
    16'h1,
    16'hffeb,
    16'h19,
    16'hfff5,
    16'hffe7,
    16'ha,
    16'hfff1,
    16'ha,
    16'h18,
    16'h7,
    16'hfffd,
    16'hffff,
    16'hfff1,
    16'hfff7,
    16'hffe4,
    16'hfff0,
    16'ha,
    16'h9,
    16'hffdd,
    16'hc,
    16'hc,
    16'hfff9,
    16'hfff3,
    16'hffe8,
    16'hffd7,
    16'h20,
    16'h12,
    16'h11,
    16'hffec,
    16'h6,
    16'h1,
    16'hfffd,
    16'h9,
    16'hfff2,
    16'ha,
    16'hfffa,
    16'hffe6,
    16'hfff8,
    16'h17,
    16'h7,
    16'h1a,
    16'hc,
    16'hffef,
    16'hffe7,
    16'h2,
    16'hfff3,
    16'hfff0,
    16'hffe7,
    16'hffcc,
    16'hfff7,
    16'hd,
    16'hffed,
    16'hffee,
    16'hfff5,
    16'h9,
    16'hffdf,
    16'hffff,
    16'hfff5,
    16'hffe9,
    16'h1d,
    16'h0,
    16'hffd9,
    16'hffe5,
    16'hb,
    16'h7,
    16'hfff5,
    16'hfff5,
    16'h29,
    16'h30,
    16'h6,
    16'h2,
    16'hffde,
    16'hfffe,
    16'h22,
    16'ha,
    16'h16,
    16'hffe8,
    16'hffe2,
    16'h2,
    16'hffee,
    16'hffff,
    16'hfffb,
    16'hffe1,
    16'hfff2,
    16'hffe1,
    16'hffec,
    16'hffe5,
    16'hfff0,
    16'hffd3,
    16'hffe2,
    16'hffef,
    16'hfff5,
    16'hfff7,
    16'h14,
    16'hfff8,
    16'hffea,
    16'hfff3,
    16'h32,
    16'h19,
    16'h9,
    16'hffd8,
    16'hffd3,
    16'h3,
    16'hffea,
    16'hfff2,
    16'h0,
    16'hfff7,
    16'hffdb,
    16'hffc8,
    16'hffe5,
    16'hfffd,
    16'h6,
    16'hfff8,
    16'h1,
    16'hfffb,
    16'h17,
    16'hffec,
    16'h9,
    16'hfff0,
    16'hfff8,
    16'hfffe,
    16'hfffc,
    16'hfff8,
    16'h26,
    16'h14,
    16'h3,
    16'hffcc,
    16'hfffc,
    16'h1d,
    16'hfff8,
    16'hf,
    16'h1d,
    16'ha,
    16'h5,
    16'h2f,
    16'h6,
    16'hffcb,
    16'hffd4,
    16'hffe9,
    16'hffe7,
    16'hfffc,
    16'hfff4,
    16'h10,
    16'h20,
    16'h0,
    16'hffe7,
    16'hfffb,
    16'hfff8,
    16'hfff7,
    16'hfff9,
    16'hc,
    16'hd,
    16'hfff7,
    16'hfff2,
    16'hffda,
    16'hffea,
    16'hffc8,
    16'hffe8,
    16'hfffb,
    16'h9,
    16'hffec,
    16'h1,
    16'hfffa,
    16'h4,
    16'hfffd,
    16'hfffb,
    16'h1b,
    16'h14,
    16'hffff,
    16'h0,
    16'hfff8,
    16'hfff2,
    16'h19,
    16'hfff7,
    16'h2,
    16'hfff9,
    16'hffef,
    16'hffed,
    16'hfff2,
    16'hfffa,
    16'he,
    16'h2,
    16'hffe5,
    16'he,
    16'hfff3,
    16'hffef,
    16'hffef,
    16'hfffb,
    16'h10,
    16'hffe7,
    16'hffe8,
    16'hffe4,
    16'he,
    16'h27,
    16'hc,
    16'hffeb,
    16'hf,
    16'h0,
    16'h22,
    16'h1e,
    16'h6,
    16'h15,
    16'h24,
    16'hfffc,
    16'h3d,
    16'h1a,
    16'h18,
    16'hffe5,
    16'hffd5,
    16'hffdd,
    16'hffdc,
    16'hfff6,
    16'h19,
    16'h12,
    16'hfffa,
    16'hffe5,
    16'hfff6,
    16'h30,
    16'hffee,
    16'h15,
    16'h7,
    16'hffc3,
    16'hffc2,
    16'hffcc,
    16'hffe7,
    16'hfff5,
    16'hffe6,
    16'h14,
    16'hfffd,
    16'hfff1,
    16'hffde,
    16'hffed,
    16'ha,
    16'h8,
    16'h5,
    16'h2c,
    16'h2,
    16'he,
    16'h7,
    16'hffe8,
    16'h6,
    16'h14,
    16'hffdb,
    16'h1e,
    16'hfff5,
    16'hffce,
    16'hc,
    16'hffd8,
    16'hb,
    16'hffe6,
    16'hffd8,
    16'h1f,
    16'h10,
    16'h1a,
    16'h11,
    16'he,
    16'hffe3,
    16'hffc3,
    16'hfff8,
    16'h35,
    16'h3,
    16'hffe4,
    16'hfff9,
    16'h2c,
    16'he,
    16'h17,
    16'h11,
    16'h3,
    16'hffeb,
    16'hffee,
    16'h2,
    16'h2,
    16'hffce,
    16'hfff1,
    16'he,
    16'hfff3,
    16'hc,
    16'hffee,
    16'hfffc,
    16'h5,
    16'h2,
    16'hb,
    16'h5,
    16'h2,
    16'hffdd,
    16'hfff2,
    16'hffef,
    16'h4,
    16'hfff9,
    16'hffe1,
    16'hffff,
    16'hffed,
    16'hffdb,
    16'h27,
    16'h9,
    16'hffe5,
    16'hffdb,
    16'hc,
    16'he,
    16'h1a,
    16'hfffc,
    16'h13,
    16'hffd3,
    16'h2,
    16'hfff5,
    16'h16,
    16'hfffa,
    16'hffff,
    16'hfffd,
    16'hffe8,
    16'h7,
    16'h1,
    16'hffff,
    16'hffc8,
    16'hffd8,
    16'h5,
    16'hffec,
    16'h6,
    16'hfffa,
    16'hffd8,
    16'hffca,
    16'h7,
    16'hffe3,
    16'hffe7,
    16'hffdc,
    16'hfffc,
    16'hf,
    16'hffe4,
    16'hfffd,
    16'h3,
    16'h18,
    16'hffe3,
    16'hffe2,
    16'ha,
    16'h25,
    16'h2d,
    16'ha,
    16'h1d,
    16'hfffe,
    16'hfffd,
    16'h24,
    16'hfff7,
    16'h15,
    16'h48,
    16'h13,
    16'hfff4,
    16'hfffc,
    16'hfffa,
    16'hffd3,
    16'hffd8,
    16'hffed,
    16'hffeb,
    16'hffe2,
    16'hfff1,
    16'hffe2,
    16'hffe6,
    16'hd,
    16'h17,
    16'h37,
    16'h30,
    16'h9,
    16'h28,
    16'h4,
    16'h16,
    16'hfff4,
    16'h6,
    16'h12,
    16'hfff4,
    16'h10,
    16'h5,
    16'hffe4,
    16'hfffe,
    16'hffec,
    16'hfffa,
    16'hfff3,
    16'hfff6,
    16'h12,
    16'hffff,
    16'hffed,
    16'hfff5,
    16'h0,
    16'hffe7,
    16'hffe2,
    16'hffe9,
    16'h11,
    16'hfffc,
    16'hffef,
    16'hffe6,
    16'hffe6,
    16'hffe3,
    16'hfffc,
    16'hffe8,
    16'hfff5,
    16'h7,
    16'hffeb,
    16'hffee,
    16'hfffd,
    16'hffe9,
    16'hfff1,
    16'hffe7,
    16'hfffa,
    16'h1e,
    16'h5d,
    16'h21,
    16'hffea,
    16'h1b,
    16'h3,
    16'hffff,
    16'hfff0,
    16'h23,
    16'he,
    16'he,
    16'h12,
    16'hfff0,
    16'hfffe,
    16'hfffb,
    16'hfff8,
    16'hfffd,
    16'hffec,
    16'hc,
    16'h6,
    16'hffde,
    16'hffdb,
    16'hffe3,
    16'hfff2,
    16'hffeb,
    16'hffe1,
    16'hfffa,
    16'hb,
    16'hfff7,
    16'hfffc,
    16'h6,
    16'h6,
    16'h2f,
    16'h2f,
    16'h13,
    16'h4,
    16'h2,
    16'h7,
    16'hffde,
    16'h2,
    16'h21,
    16'h2d,
    16'h2e,
    16'h30,
    16'hffec,
    16'hfff4,
    16'hffdb,
    16'hffb6,
    16'hffef,
    16'h14,
    16'hfff5,
    16'hffe9,
    16'hffd8,
    16'hffff,
    16'h17,
    16'hffeb,
    16'ha,
    16'hfff8,
    16'h9,
    16'h2b,
    16'h21,
    16'h15,
    16'h0,
    16'hfff6,
    16'h1,
    16'h7,
    16'hffe4,
    16'hffe6,
    16'h2,
    16'h6,
    16'h8,
    16'hffe7,
    16'hfff0,
    16'h9,
    16'h16,
    16'hfff0,
    16'h18,
    16'hffff,
    16'hfff7,
    16'hfff4,
    16'h1,
    16'hffec,
    16'hffee,
    16'hffea,
    16'h4,
    16'h12,
    16'h14,
    16'hb,
    16'hffcb,
    16'hffd0,
    16'hffe6,
    16'hffe0,
    16'h8,
    16'hfff4,
    16'hc,
    16'hfff0,
    16'h1,
    16'hf,
    16'hffed,
    16'h10,
    16'hf,
    16'he,
    16'hc,
    16'hfffc,
    16'h3,
    16'hfff4,
    16'h15,
    16'h18,
    16'hfffb,
    16'hffd4,
    16'hffef,
    16'hfffc,
    16'hffdf,
    16'hfff2,
    16'hd,
    16'h21,
    16'hc,
    16'h0,
    16'hfffe,
    16'h1d,
    16'h2c,
    16'h9,
    16'hb,
    16'h15,
    16'ha,
    16'h9,
    16'hffda,
    16'hfffe,
    16'h10,
    16'h9,
    16'hffdf,
    16'hfff5,
    16'hfff2,
    16'h11,
    16'hb,
    16'hfff7,
    16'hd,
    16'h4,
    16'hfffa,
    16'h2,
    16'hffe2,
    16'h1,
    16'hc,
    16'hffe9,
    16'hfffe,
    16'h3,
    16'h20,
    16'hfff9,
    16'h6,
    16'hffd4,
    16'hffdd,
    16'h9,
    16'hfff9,
    16'h1d,
    16'hfff7,
    16'hffd8,
    16'hfff5,
    16'hfff2,
    16'hffd8,
    16'hffed,
    16'h6,
    16'hfff5,
    16'h24,
    16'hffe8,
    16'hffff,
    16'h15,
    16'hfff7,
    16'h8,
    16'h17,
    16'hfff5,
    16'he,
    16'h10,
    16'hfff6,
    16'hfff4,
    16'hffd8,
    16'hfffa,
    16'hfffb,
    16'h2,
    16'ha,
    16'h16,
    16'hfff9,
    16'hffe8,
    16'h15,
    16'hffe5,
    16'hfffc,
    16'hffef,
    16'hfffb,
    16'hfffd,
    16'hfff8,
    16'hffeb,
    16'hfffc,
    16'hfff5,
    16'hfff3,
    16'hffe0,
    16'hffe2,
    16'hffe4,
    16'h6,
    16'h9,
    16'h9,
    16'hffee,
    16'hffe9,
    16'hb,
    16'h13,
    16'hfff0,
    16'h12,
    16'hd,
    16'hffee,
    16'h17,
    16'h7,
    16'h15,
    16'h6,
    16'h17,
    16'hffea,
    16'h11,
    16'h7,
    16'h10,
    16'hfff3,
    16'hffd0,
    16'hffe0,
    16'hfffc,
    16'h14,
    16'hffda,
    16'hffc8,
    16'hffd7,
    16'ha,
    16'h3,
    16'h0,
    16'hd,
    16'hffcc,
    16'h27,
    16'h41,
    16'h3d,
    16'h1a,
    16'h8,
    16'hffbc,
    16'h0,
    16'h2d,
    16'h7,
    16'hb,
    16'h1,
    16'hffdd,
    16'hb,
    16'hfff9,
    16'hb,
    16'hfff1,
    16'hfffd,
    16'h3,
    16'h24,
    16'h1b,
    16'h17,
    16'hfff6,
    16'h9,
    16'h1,
    16'h1d,
    16'h4,
    16'hffeb,
    16'h10,
    16'h6,
    16'hfff8,
    16'hffb8,
    16'hfffc,
    16'h14,
    16'h12,
    16'hffd5,
    16'hffe1,
    16'hfffb,
    16'hffe9,
    16'hffe6,
    16'hfffb,
    16'hfff3,
    16'hfff9,
    16'hffeb,
    16'hffe5,
    16'hfffa,
    16'h7,
    16'h19,
    16'h1d,
    16'h14,
    16'hffff,
    16'hb,
    16'hffec,
    16'h9,
    16'hfff9,
    16'hfff2,
    16'hffe1,
    16'hffec,
    16'hffec,
    16'h6,
    16'hf,
    16'hffec,
    16'ha,
    16'hfffb,
    16'ha,
    16'hffe0,
    16'h1f,
    16'h23,
    16'h1f,
    16'hffe8,
    16'ha,
    16'hfff5,
    16'hffff,
    16'hfffe,
    16'hfffd,
    16'hfff1,
    16'h17,
    16'h12,
    16'h33,
    16'h25,
    16'hc,
    16'hffee,
    16'hfff9,
    16'h16,
    16'h1a,
    16'hffe8,
    16'hffd9,
    16'hffee,
    16'h1,
    16'hfffa,
    16'hffc3,
    16'hffcc,
    16'hffe6,
    16'ha
  };
  // logic signed [15:0] threshold [0:OC-1] = {-16'd31, -16'd73, -16'd16, -16'd33, -16'd13, -16'd3, -16'd1543, -16'd4, -16'd8, -16'd14};
  // logic [CONV1_IMG_OUT_SIZE*CONV1_IMG_OUT_SIZE-1:0] conv1_img_out [0:CONV1_OC-1];
  logic [POOL1_IMG_OUT_SIZE*POOL1_IMG_OUT_SIZE-1:0] pool1_img_out[0:CONV1_OC-1];
  // logic [CONV2_IMG_OUT_SIZE*CONV2_IMG_OUT_SIZE-1:0] conv2_img_out [0:CONV2_OC-1];
  logic [POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE-1:0] pool2_img_out[0:CONV2_OC-1];
  logic [FC_IC-1:0] fc_in;
  logic signed [15:0] fc_out[0:FC_OC-1];
  logic conv1_data_ready;
  // logic pool1_data_ready;
  logic conv2_data_ready;
  // logic pool2_data_ready;
  logic fc_data_ready;

  Conv2d_MaxPool2d #(
      .IC(CONV1_IC),
      .OC(CONV1_OC),
      .CONV_IMG_IN_SIZE(CONV1_IMG_IN_SIZE)
  ) conv_pool1 (
      .clk(clk),
      .data_in_ready(data_in_ready),
      .img_in(conv1_img_in),
      .weights(conv1_weights),
      .img_out(pool1_img_out),
      .data_out_ready(conv1_data_ready)
  );

  Conv2d_MaxPool2d #(
      .IC(CONV1_OC),
      .OC(CONV2_OC),
      .CONV_IMG_IN_SIZE(POOL1_IMG_OUT_SIZE)
  ) conv_pool2 (
      .clk(clk),
      .data_in_ready(conv1_data_ready),
      .img_in(pool1_img_out),
      .weights(conv2_weights),
      .img_out(pool2_img_out),
      .data_out_ready(conv2_data_ready)
  );

  genvar conv2_oc;
  generate
    for (conv2_oc = 0; conv2_oc < CONV2_OC; conv2_oc = conv2_oc + 1) begin
      assign fc_in[conv2_oc*POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE +: POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE] = pool2_img_out[conv2_oc];
    end
  endgenerate


  FC #(
      .IC(FC_IC),
      .OC(FC_OC)
  ) fc (
      .clk(clk),
      .data_in_ready(conv2_data_ready),
      .in(fc_in),
      .weights(fc_weights),
      .out(fc_out),
      .data_out_ready(fc_data_ready)
  );

  Comparator #(
      .IC(FC_OC)
  ) compare (
      .clk(clk),
      .data_in_ready(fc_data_ready),
      .in(fc_out),
      .out(result),
      .data_out_ready(data_out_ready)
  );

  // wire _unused_ok = &{result};

endmodule
