`include "Conv2d.sv"
`include "MaxPool2d.sv"

module bnn_top (
    // input logic [CONV1_IMG_IN_SIZE*CONV1_IMG_IN_SIZE-1:0] img_in [0:CONV1_IC-1]
    input logic clk,
    input logic data_in_ready,
    output logic [OUTPUT_BIT-1:0] result,
    output logic data_out_ready
);
    parameter int CONV1_IC = 1;
    parameter int CONV1_OC = 10;
    parameter int CONV2_OC = 8;
    parameter int FC_IC= POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE*CONV2_OC;
    parameter int FC_OC = 10;                   // num classes
    parameter int CONV1_IMG_IN_SIZE = 30;
    parameter int CONV1_IMG_OUT_SIZE = CONV1_IMG_IN_SIZE-2;
    parameter int POOL1_IMG_OUT_SIZE = CONV1_IMG_OUT_SIZE/2;
    parameter int CONV2_IMG_OUT_SIZE = POOL1_IMG_OUT_SIZE-2;
    parameter int POOL2_IMG_OUT_SIZE = CONV2_IMG_OUT_SIZE/2;
    parameter int OUTPUT_BIT = $clog2(FC_OC+1); // num of bits to enumerate each class

    logic [CONV1_IMG_IN_SIZE*CONV1_IMG_IN_SIZE-1:0] conv1_img_in [0:CONV1_IC-1] = {900'h7c000003fc00001e70000070000001800000070000001ff000001fe0000001800000060000081800003ff00000ffc0000000000000000000000000000000000000000000000000000000000000000000000};
    // assign conv1_img_in = img_in;
    logic [CONV1_IC*9-1:0] conv1_weights [0:CONV1_OC-1] = {9'hb5, 9'h180, 9'h1ef, 9'h3c, 9'h108, 9'hdb, 9'hdf, 9'h120, 9'h1e9, 9'h5f};
    logic [CONV1_OC*9-1:0] conv2_weights [0:CONV2_OC-1] = {90'hb5b844a62f6db494cd83fa, 90'hbf8800fff4800007b4056e, 90'h9440867301210005b60924, 90'h2b209cb22cbf7fcfc16a769, 90'hafd05355b11c000f7591c6, 90'h7d80d18fc0f22200140026, 90'h23962017fef20823ffe4fbc, 90'h3baed0113c928200791332c};
    logic signed [15:0] fc_weights [0:FC_IC*FC_OC-1] = {16'hffde, 16'hc, 16'h20, 16'h20, 16'ha, 16'hffd0, 16'hfffc, 16'h9, 16'h1c, 16'hb, 16'hfffa, 16'hffeb, 16'h25, 16'h34, 16'h2a, 16'h1d, 16'h3c, 16'h47, 16'hf, 16'hfffc, 16'h2d, 16'h35, 16'h77, 16'h4d, 16'hfffc, 16'hfff2, 16'h1d, 16'h3a, 16'h3d, 16'h24, 16'hfff2, 16'h11, 16'hfffc, 16'hffed, 16'h13, 16'hfff2, 16'hfff5, 16'hffd5, 16'hffd3, 16'hffff, 16'hffe5, 16'hffe1, 16'hffee, 16'hffc6, 16'hffcb, 16'hffa7, 16'hff98, 16'h1b, 16'hffd6, 16'hffca, 16'hff5a, 16'hff5a, 16'hff3d, 16'hffea, 16'hffe5, 16'hffb9, 16'hff4f, 16'hff40, 16'hff3d, 16'hffb7, 16'hfff3, 16'hd, 16'hffb8, 16'hffab, 16'hffa4, 16'hfffe, 16'hfff1, 16'h15, 16'h5, 16'h1c, 16'h18, 16'h6, 16'hffd8, 16'hffc5, 16'hffde, 16'hffe7, 16'h7, 16'h1, 16'hffcd, 16'hffd4, 16'h6, 16'h30, 16'h20, 16'h10, 16'hffee, 16'hd, 16'h76, 16'h8b, 16'h5b, 16'h9, 16'h42, 16'h59, 16'hb0, 16'h7a, 16'h35, 16'hfff1, 16'h39, 16'h44, 16'h5e, 16'h3a, 16'hfff2, 16'hffef, 16'hffff, 16'h14, 16'h7, 16'hffe7, 16'hffb5, 16'hffd5, 16'h1c, 16'h3c, 16'h2e, 16'hffef, 16'h1, 16'h5, 16'hf, 16'hfff1, 16'hffe9, 16'hfff6, 16'h37, 16'hc, 16'h2d, 16'hffe5, 16'hffcc, 16'hffed, 16'hfff0, 16'hffd9, 16'hf, 16'hffc6, 16'hffbf, 16'hffdf, 16'hfff6, 16'hffd0, 16'h3b, 16'hffec, 16'h14, 16'hffe5, 16'hffe0, 16'hffe1, 16'h14, 16'hffed, 16'h2b, 16'hf, 16'h6, 16'hfffc, 16'hfffe, 16'hffe6, 16'hffda, 16'h1c, 16'h16, 16'h6, 16'hffef, 16'hffe8, 16'h1, 16'h14, 16'h3f, 16'h4a, 16'h21, 16'ha, 16'h8, 16'h0, 16'h2a, 16'h43, 16'hffd1, 16'hffdf, 16'hfff4, 16'hfff5, 16'h2, 16'h12, 16'hffba, 16'hffee, 16'h8, 16'hffeb, 16'hffec, 16'hffec, 16'hffce, 16'hfff8, 16'h4, 16'hffe1, 16'hffef, 16'hffe2, 16'hffd9, 16'hfff1, 16'hffff, 16'hfff0, 16'hffeb, 16'hfff3, 16'hffd3, 16'hffb1, 16'hffe5, 16'h4f, 16'h54, 16'h16, 16'hffdb, 16'hff9a, 16'hffbf, 16'hfff2, 16'h17, 16'h5, 16'hfffd, 16'hffce, 16'hffd3, 16'hffd4, 16'hffe2, 16'he, 16'hd, 16'hfff9, 16'hffea, 16'hffdf, 16'hffda, 16'hfff1, 16'he, 16'h17, 16'hfffe, 16'hfffa, 16'hffef, 16'hfff9, 16'h3, 16'hffc6, 16'h32, 16'h79, 16'h3b, 16'h3, 16'hffd8, 16'h39, 16'h21, 16'h34, 16'h3a, 16'h3f, 16'hffee, 16'h7f, 16'h7b, 16'h49, 16'h32, 16'h43, 16'h41, 16'h9a, 16'h66, 16'h1e, 16'h16, 16'h43, 16'h4d, 16'h69, 16'h25, 16'h13, 16'h2e, 16'h28, 16'hffd9, 16'h38, 16'h17, 16'h1f, 16'h41, 16'hd, 16'hffe2, 16'hb, 16'he, 16'h21, 16'h54, 16'h1a, 16'h8, 16'hfffd, 16'hfffc, 16'h1b, 16'h7a, 16'h65, 16'hffcf, 16'hfff6, 16'h1d, 16'h37, 16'h4f, 16'h40, 16'hfff2, 16'hd, 16'h3b, 16'h3d, 16'h19, 16'h16, 16'hffcb, 16'h16, 16'h3a, 16'h34, 16'hfffa, 16'h7, 16'h5, 16'h2, 16'h22, 16'h40, 16'ha, 16'hffef, 16'hf, 16'hff9b, 16'hffc3, 16'hfffc, 16'hffa2, 16'h0, 16'hffda, 16'hff91, 16'hffca, 16'hffe1, 16'hff87, 16'hffb4, 16'hffbd, 16'hffaa, 16'hff79, 16'hff7f, 16'hff85, 16'hffa4, 16'hffdd, 16'hff94, 16'hffa2, 16'hff9c, 16'hff76, 16'hffa5, 16'hffcd, 16'hffd4, 16'hffcd, 16'hffce, 16'hffa8, 16'hffc9, 16'hfff3, 16'hfff8, 16'hffed, 16'hffdc, 16'hffd5, 16'hffc8, 16'h6, 16'h33, 16'hffea, 16'h3, 16'hfff4, 16'h40, 16'h1e, 16'h17, 16'hc, 16'hfffa, 16'h20, 16'h4, 16'h39, 16'hfff4, 16'hffe6, 16'h32, 16'h1c, 16'hfff2, 16'h2e, 16'hffd6, 16'hff9e, 16'hffde, 16'hffff, 16'h1, 16'h2d, 16'h0, 16'hffa2, 16'hffce, 16'hffe6, 16'h23, 16'h3e, 16'hfff5, 16'hffeb, 16'hffd7, 16'hffed, 16'h38, 16'h1b, 16'h23, 16'h15, 16'h2c, 16'hd, 16'hb, 16'h29, 16'hffeb, 16'hc, 16'h1f, 16'h14, 16'hfff6, 16'hffe7, 16'hffd9, 16'h1f, 16'hb, 16'h7, 16'h2, 16'h2, 16'hfff5, 16'h27, 16'h35, 16'hfff4, 16'h15, 16'hfff6, 16'h1a, 16'h34, 16'h35, 16'h0, 16'h20, 16'h4, 16'h29, 16'h24, 16'h37, 16'h14, 16'ha, 16'hffe1, 16'hfff2, 16'hffe7, 16'hfffe, 16'hffd3, 16'hffff, 16'hfffe, 16'hfffa, 16'hffe9, 16'hff9e, 16'hfff4, 16'hffda, 16'hfff3, 16'h2, 16'hffd0, 16'hffb2, 16'hffd9, 16'hffd2, 16'hffba, 16'hffe6, 16'hffc5, 16'hffd6, 16'hffd7, 16'hffc3, 16'hffd2, 16'hffeb, 16'hffd3, 16'hfff6, 16'hfff5, 16'hffbd, 16'hfffe, 16'hffe0, 16'hffe9, 16'hffec, 16'hfffb, 16'hffd5, 16'h8, 16'hffc9, 16'hffc9, 16'hfff6, 16'hffd0, 16'hffca, 16'h30, 16'hffb0, 16'hff8c, 16'hffc6, 16'hffc3, 16'hffc5, 16'hffe8, 16'hffd8, 16'hffb4, 16'hffa3, 16'hffc9, 16'hffc4, 16'h22, 16'hfffa, 16'hffb6, 16'hffc5, 16'hffc1, 16'hffd6, 16'h21, 16'hfff0, 16'hffe2, 16'hffdf, 16'hffe4, 16'hffe8, 16'h3a, 16'hfffa, 16'hfffe, 16'h7, 16'hfff9, 16'h8, 16'h41, 16'h1e, 16'h27, 16'h39, 16'h42, 16'h48, 16'h11, 16'hffdb, 16'hffde, 16'hfffe, 16'hfff3, 16'h1b, 16'hffe7, 16'hffdc, 16'h6, 16'hffe6, 16'hffd1, 16'h21, 16'hffd2, 16'hffbb, 16'hffdc, 16'hffc3, 16'hffe7, 16'h11, 16'hffc7, 16'hffe2, 16'hffc1, 16'hffcd, 16'hffe3, 16'hfff8, 16'hffe2, 16'hd, 16'hfff9, 16'h8, 16'hfff5, 16'h12, 16'h3c, 16'hfff7, 16'hff9f, 16'hff77, 16'hffa6, 16'h14, 16'h14, 16'h1, 16'hffc4, 16'hff9b, 16'hffb3, 16'hffe4, 16'h0, 16'hffd8, 16'hffa6, 16'hff9d, 16'hff95, 16'hffbd, 16'h23, 16'hffe3, 16'hffc2, 16'hffa6, 16'hffa8, 16'hffc8, 16'h2b, 16'hffe8, 16'hffc2, 16'hff9e, 16'hff9a, 16'hffd4, 16'h2e, 16'hffdf, 16'hff8f, 16'hff74, 16'hffc6, 16'hffcf, 16'h7, 16'h3, 16'h1f, 16'hffe9, 16'h7, 16'hffdf, 16'hf, 16'h2e, 16'hffea, 16'h2c, 16'h4f, 16'h11, 16'h2c, 16'h13, 16'hffb9, 16'hfff8, 16'h2a, 16'h4, 16'h2f, 16'hfff4, 16'hffd1, 16'hfff0, 16'h33, 16'h2a, 16'h3d, 16'hfffa, 16'hffc3, 16'hffd4, 16'h4, 16'h1e, 16'h29, 16'h2, 16'hffed, 16'hffe7, 16'hfff4, 16'hfffc, 16'h6, 16'h15, 16'h10, 16'hffca, 16'hffb7, 16'hffdd, 16'hffbb, 16'h32, 16'hf, 16'hff8b, 16'hffaa, 16'hffe4, 16'hd, 16'h16, 16'hffec, 16'hffe8, 16'hffe5, 16'h11, 16'h64, 16'h85, 16'h60, 16'h3f, 16'h51, 16'h4e, 16'h4b, 16'h88, 16'h5f, 16'hffd7, 16'hfffa, 16'h17, 16'h18, 16'h38, 16'hffe6, 16'hffb6, 16'hffe2, 16'h17, 16'hffe7, 16'h15, 16'hffff, 16'hffd7, 16'hffd0, 16'hd, 16'hffeb, 16'hffba, 16'hff8b, 16'hff5f, 16'hff63, 16'hfff5, 16'h14, 16'hffd4, 16'hffc1, 16'hffa1, 16'hff7c, 16'hffd5, 16'h19, 16'hffd6, 16'h17, 16'hf, 16'hffee, 16'hfffd, 16'hc, 16'hffd1, 16'h55, 16'h78, 16'h43, 16'h2d, 16'h12, 16'hfffd, 16'h14, 16'h5c, 16'h26, 16'h14, 16'h6, 16'h0, 16'h21, 16'h4b, 16'h30, 16'h25, 16'h0, 16'hffed, 16'hffd3, 16'h4a, 16'h34, 16'h15, 16'hffa7, 16'hffcb, 16'hffab, 16'h6, 16'h17, 16'h16, 16'hffd2, 16'hffc6, 16'hffad, 16'hffd3, 16'hfffd, 16'hfffb, 16'hffec, 16'hffc5, 16'hffae, 16'hffa6, 16'hffcf, 16'hfff1, 16'he, 16'hffe9, 16'hffd0, 16'hffb6, 16'hffe9, 16'h15, 16'hfff6, 16'hfffb, 16'h3, 16'h1e, 16'hfffb, 16'hfff5, 16'h2a, 16'h30, 16'h52, 16'h24, 16'h24, 16'h21, 16'h10, 16'h3e, 16'h4e, 16'h1, 16'hffe3, 16'h10, 16'hfff2, 16'h65, 16'h1d, 16'hfff6, 16'hffdf, 16'hfff7, 16'hfffa, 16'h2a, 16'h2, 16'hffec, 16'h3, 16'h2e, 16'hf, 16'hfffb, 16'hfff9, 16'h22, 16'ha, 16'h13, 16'hfff5, 16'h0, 16'h2d, 16'h16, 16'hffdf, 16'hffc8, 16'hffef, 16'h20, 16'hfff1, 16'hffc5, 16'hffdb, 16'hffe0, 16'h67, 16'h69, 16'hffb7, 16'hffa6, 16'hfffd, 16'h3, 16'h52, 16'h20, 16'hff95, 16'hffa8, 16'hffe6, 16'hffef, 16'h40, 16'h19, 16'hffc1, 16'hffbe, 16'hfff7, 16'hfffc, 16'hfff8, 16'hffbc, 16'hff94, 16'hff9f, 16'hffee, 16'h25, 16'hfff0, 16'hfff5, 16'h2, 16'hffc8, 16'hfff2, 16'hffd7, 16'hfff8, 16'h79, 16'ha3, 16'h6d, 16'h2f, 16'hfffe, 16'hc, 16'h54, 16'h76, 16'h42, 16'h1c, 16'hffde, 16'h44, 16'h69, 16'h55, 16'h5e, 16'h6f, 16'h71, 16'h43, 16'h2e, 16'ha, 16'h32, 16'h42, 16'h59, 16'h24, 16'h19, 16'hfffd, 16'h7, 16'h31, 16'h49, 16'h11, 16'hffd0, 16'hfffe, 16'h25, 16'hfff4, 16'hffde, 16'hfff9, 16'hff70, 16'hffb8, 16'hfffc, 16'hffff, 16'hfff1, 16'hffc7, 16'hff65, 16'hff93, 16'hfff9, 16'hfffc, 16'h1, 16'hffa5, 16'hffc0, 16'hffde, 16'h16, 16'h25, 16'h4, 16'hffc5, 16'hfff7, 16'hffe3, 16'h38, 16'ha, 16'h16, 16'hc, 16'hc, 16'hffdd, 16'hfffd, 16'h2d, 16'h24, 16'hfff9, 16'hfffa, 16'hffed, 16'h23, 16'h20, 16'h20, 16'hffdc, 16'h19, 16'hffd3, 16'h14, 16'h32, 16'h21, 16'hc, 16'h38, 16'h13, 16'hffef, 16'hffd8, 16'hffc4, 16'hfffe, 16'h77, 16'h2f, 16'hffe8, 16'hffc5, 16'hffa4, 16'hd, 16'h44, 16'h3b, 16'h2d, 16'hffdd, 16'hffa6, 16'h18, 16'h3e, 16'h3b, 16'h4d, 16'h2, 16'hfff1, 16'h11, 16'h50, 16'hfff6, 16'hffec, 16'hffe0, 16'hffdc, 16'hffbd, 16'h1a, 16'h20, 16'hfff0, 16'hffe9, 16'hffff, 16'hffd1, 16'hffe1, 16'hff9f, 16'h0, 16'hffef, 16'hfff7, 16'h4d, 16'h52, 16'h3e, 16'h50, 16'hfff7, 16'hffca, 16'h47, 16'h7e, 16'h90, 16'h46, 16'hffdc, 16'hffcd, 16'h30, 16'h46, 16'h2e, 16'h22, 16'hffe4, 16'hffcb, 16'h28, 16'hffef, 16'h1, 16'h4, 16'h25, 16'h10, 16'hffef, 16'hfffd, 16'hfff8, 16'h25, 16'h6e, 16'h10, 16'hfff0, 16'hfff5, 16'hffff, 16'h44, 16'h84, 16'h21, 16'h1a, 16'hffe3, 16'hff86, 16'hffd5, 16'h1f, 16'h17, 16'h5, 16'hffc7, 16'hff46, 16'hff53, 16'hffa9, 16'h11, 16'ha, 16'h2, 16'hff9d, 16'hffae, 16'hffe7, 16'hfff7, 16'h9, 16'hfff7, 16'h1b, 16'hffff, 16'h2a, 16'h1e, 16'h28, 16'hffd1, 16'hffd4, 16'hffdd, 16'h18, 16'h8, 16'hffcc, 16'hffcf, 16'hffd2, 16'hffc4, 16'hfff1, 16'hfffc, 16'hffd8, 16'hffc7, 16'hffe3, 16'hffdc, 16'hffd1, 16'hffd5, 16'h17, 16'hfff2, 16'hfffa, 16'hffdb, 16'hffe1, 16'hffe3, 16'h1f, 16'h11, 16'hfff3, 16'hffdf, 16'hffe4, 16'hfffb, 16'hffd9, 16'hb, 16'hffd3, 16'hfff5, 16'hffe9, 16'hffd2, 16'hffd9, 16'hf, 16'h65, 16'h25, 16'hfff9, 16'h9, 16'hfff9, 16'h2f, 16'h73, 16'h36, 16'h7, 16'h15, 16'h6, 16'h3a, 16'h54, 16'h33, 16'hfffb, 16'hfff8, 16'hffe2, 16'h2f, 16'h32, 16'h15, 16'hfff3, 16'h8, 16'hfff9, 16'hfffd, 16'h2, 16'hffed, 16'h6, 16'hffe4, 16'he, 16'h28, 16'h19, 16'hfff3, 16'hfff8, 16'h4, 16'hffff, 16'hfffc, 16'hffec, 16'hfff2, 16'he, 16'h26, 16'hffff, 16'h33, 16'h13, 16'h3, 16'hfffa, 16'h3, 16'h45, 16'h8a, 16'h66, 16'h2a, 16'hffec, 16'hffd5, 16'h54, 16'h9d, 16'ha1, 16'h2d, 16'hffe4, 16'hffd7, 16'hffed, 16'hd, 16'he, 16'hffe9, 16'hffd1, 16'hffd5, 16'h2, 16'h26, 16'h9, 16'hffe5, 16'hffe5, 16'h1b, 16'hffeb, 16'h76, 16'h4d, 16'hffea, 16'hffc5, 16'hffff, 16'hfff0, 16'h37, 16'h4d, 16'hffec, 16'hffe6, 16'hfff5, 16'h9, 16'h1, 16'h3b, 16'h34, 16'hfff7, 16'hffb7, 16'h42, 16'h49, 16'h60, 16'h2a, 16'hffd7, 16'hffad, 16'h2a, 16'h2b, 16'h2c, 16'h8, 16'hffe8, 16'hfff1, 16'hffee, 16'hffe3, 16'hd, 16'h28, 16'hd, 16'h27, 16'hfff1, 16'hff81, 16'hffd1, 16'h5b, 16'h32, 16'h4e, 16'h7, 16'hff21, 16'hff5e, 16'hffeb, 16'h8, 16'h3a, 16'hffdd, 16'hff57, 16'hff73, 16'hffbb, 16'hfff4, 16'hc, 16'hffc5, 16'hffb7, 16'hffc0, 16'h9, 16'h24, 16'h3, 16'h8, 16'hf, 16'h36, 16'h30, 16'h33, 16'h5, 16'h18, 16'hffec, 16'h10, 16'hffdf, 16'h37, 16'h1c, 16'hf, 16'h2f, 16'hfff0, 16'hffe9, 16'h17, 16'h15, 16'h2f, 16'hfff6, 16'hffd6, 16'hffd0, 16'hfffb, 16'h18, 16'h13, 16'ha, 16'hffe9, 16'hffce, 16'hfff5, 16'hb, 16'hfff6, 16'hffe8, 16'hffea, 16'hffed, 16'hffed, 16'h1a, 16'hb, 16'h17, 16'h29, 16'h3e, 16'h1f, 16'hffe4, 16'hffd5, 16'hff8b, 16'hffbe, 16'h24, 16'h13, 16'hfffd, 16'h2c, 16'hfff5, 16'hffa7, 16'hfffd, 16'hffe1, 16'hb, 16'h79, 16'he5, 16'h46, 16'ha, 16'h1a, 16'h3f, 16'h1c, 16'h5b, 16'h38, 16'hffef, 16'h37, 16'h3b, 16'hffd9, 16'hffbd, 16'hff93, 16'hffaa, 16'hc, 16'h35, 16'hffd1, 16'hffa8, 16'hffa5, 16'hffd2, 16'hfff9, 16'hfff2, 16'hffdb, 16'h18, 16'hfff2, 16'hd, 16'h9, 16'h18, 16'hffda, 16'hffee, 16'h4d, 16'h6e, 16'h5e, 16'h24, 16'h2, 16'h34, 16'h20, 16'h3d, 16'h7, 16'h9, 16'hfff8, 16'h44, 16'h58, 16'h40, 16'h1e, 16'hffe9, 16'h0, 16'hb, 16'h79, 16'h9b, 16'h4c, 16'h15, 16'h4, 16'hffec, 16'hffeb, 16'h4, 16'h7, 16'hffe7, 16'hc, 16'h3, 16'h14, 16'hffee, 16'h33, 16'h20, 16'hffec, 16'h17, 16'h32, 16'h19, 16'h10, 16'h19, 16'hffe1, 16'hffec, 16'hffcc, 16'h1c, 16'h1a, 16'hf, 16'h6, 16'hffbf, 16'hffb8, 16'h5, 16'h11, 16'h13, 16'h4, 16'hffe1, 16'hffe7, 16'hf, 16'ha, 16'h0, 16'hffae, 16'hffd8, 16'h6, 16'h3e, 16'h34, 16'h14, 16'hffe6, 16'hfff9, 16'h11, 16'hfff3, 16'hfff1, 16'hf, 16'h14, 16'h13, 16'hff9f, 16'hffcc, 16'ha, 16'h16, 16'h1b, 16'h37, 16'hffc6, 16'hffd1, 16'hffdf, 16'h1c, 16'hffee, 16'hffdf, 16'hffc0, 16'hffea, 16'hffed, 16'h25, 16'hfffb, 16'h13, 16'h2e, 16'h3d, 16'h32, 16'h2d, 16'hfff9, 16'h22, 16'hfff1, 16'hfff6, 16'hc, 16'hfff7, 16'hffdb, 16'hffaf, 16'hff7f, 16'hffab, 16'hffe1, 16'hf, 16'h16, 16'hffee, 16'hffc4, 16'hffdb, 16'hffff, 16'h2b, 16'hfffa, 16'hffc4, 16'hffdd, 16'hffc5, 16'h3, 16'h7, 16'h7, 16'hffca, 16'hffb6, 16'hfffc, 16'h24, 16'h15, 16'hffee, 16'hffb7, 16'hffb5, 16'hffd6, 16'hfffd, 16'h3, 16'hffe3, 16'hffd7, 16'hffe1, 16'hb, 16'h6, 16'h1, 16'h16, 16'hfff1, 16'h13, 16'hfffa, 16'hffe3, 16'hffe8, 16'hffbc, 16'hff76, 16'hff54, 16'hff91, 16'hffc2, 16'h4, 16'h3b, 16'h3, 16'hffe3, 16'h1b, 16'h3d, 16'h35, 16'h5b, 16'h6b, 16'h1d, 16'he, 16'h3e, 16'h43, 16'hc, 16'hfffb, 16'hffe1, 16'h10, 16'h35, 16'h2e, 16'hfff1, 16'hffe2, 16'hffef, 16'hffec, 16'h3, 16'hfff7, 16'hffdf, 16'hffc1, 16'hff60, 16'hff9c, 16'hffbf, 16'hffe3, 16'hffe6, 16'h28, 16'hff71, 16'hff4a, 16'hffcc, 16'h41, 16'h1, 16'h6e, 16'h66, 16'h4a, 16'h21, 16'h12, 16'hfff8, 16'h14, 16'h3, 16'hffe2, 16'hfffc, 16'hfff9, 16'hffd6, 16'h10, 16'h0, 16'h16, 16'hffe4, 16'hfffc, 16'hfff7, 16'hffdf, 16'hffa7, 16'hffb3, 16'hffd9, 16'hffc5, 16'h11, 16'hffdd, 16'hffec, 16'h6, 16'h48, 16'h33, 16'h8, 16'h7, 16'h50, 16'h4e, 16'h78, 16'h47, 16'hffed, 16'h3c, 16'h4c, 16'h18, 16'h36, 16'h18, 16'hffff, 16'h0, 16'h35, 16'h10, 16'h5, 16'hffe3, 16'hb, 16'hffed, 16'h41, 16'h35, 16'hffea, 16'hffe9, 16'h3, 16'hfffb, 16'hffc3, 16'hffa9, 16'hffbd, 16'hfff1, 16'hc, 16'h26, 16'hffdd, 16'hffce, 16'h62, 16'h7b, 16'h19, 16'h1b, 16'hffe1, 16'hffc4, 16'h5c, 16'h66, 16'hffcf, 16'hffed, 16'h32, 16'h28, 16'h62, 16'h72, 16'hffc8, 16'he, 16'h18, 16'h1f, 16'h2e, 16'h2f, 16'hd, 16'h38, 16'h2e, 16'h45, 16'h26, 16'h24, 16'h1b, 16'h34, 16'h2c, 16'h29, 16'h13, 16'hfffb, 16'h11, 16'hfffa, 16'h2, 16'hffdd, 16'hffd3, 16'hfff6, 16'h26, 16'hc, 16'h2b, 16'h16, 16'hffd1, 16'hffe3, 16'hb, 16'h22, 16'hfff9, 16'hfff2, 16'hffde, 16'hffec, 16'h2a, 16'hffc9, 16'hffbc, 16'hff97, 16'hff96, 16'hffe2, 16'h26, 16'hffc4, 16'hffa6, 16'hff9f, 16'hffa9, 16'hb, 16'hffe6, 16'hffeb, 16'hffd4, 16'hffd1, 16'hffec, 16'h4, 16'h13, 16'h8, 16'h1, 16'hffc9, 16'hffc7, 16'hfff5, 16'hf, 16'h71, 16'h3d, 16'hffc7, 16'hffcc, 16'hffdf, 16'h36, 16'h66, 16'h4a, 16'hffd9, 16'hffd7, 16'hffd6, 16'ha, 16'hfffc, 16'hfff4, 16'hffd5, 16'h1, 16'hd, 16'hffdd, 16'hffc7, 16'hffc7, 16'hffc4, 16'hfff7, 16'hfffe, 16'h7, 16'hfffa, 16'hffe4, 16'hffe3, 16'hffd6, 16'hffda, 16'hfff9, 16'hffea, 16'hfffb, 16'h2, 16'hffec, 16'hffec, 16'hffe1, 16'hffca, 16'hffeb, 16'h33, 16'h1d, 16'hc, 16'h3, 16'h6, 16'hb, 16'h4f, 16'h43, 16'h3, 16'h0, 16'h22, 16'h48, 16'h3f, 16'h2e, 16'hffe9, 16'h1b, 16'h0, 16'h32, 16'he, 16'hb, 16'h9, 16'h18, 16'hf, 16'hffea, 16'hffe3, 16'hffed, 16'h8, 16'he, 16'h3c, 16'h38, 16'hfff9, 16'h21, 16'h0, 16'hffea, 16'ha, 16'h26, 16'h23, 16'h9, 16'h2, 16'hfff6, 16'hffee, 16'h47, 16'h3d, 16'h1d, 16'hfffe, 16'h36, 16'h84, 16'h72, 16'h49, 16'h21, 16'h11, 16'h18, 16'h92, 16'h80, 16'h36, 16'hfff3, 16'hffe3, 16'h2, 16'h24, 16'h1f, 16'h1, 16'hffd8, 16'hffc8, 16'hffde, 16'hfffd, 16'hfff5, 16'h5, 16'h34, 16'hffe4, 16'hfff2, 16'hffdf, 16'hfff4, 16'h73, 16'h7f, 16'h16, 16'h2a, 16'h15, 16'h3b, 16'h58, 16'h63, 16'h12, 16'hd, 16'h15, 16'h43, 16'h44, 16'h3e, 16'h19, 16'h9, 16'h34, 16'h34, 16'h39, 16'h1e, 16'h6, 16'h7, 16'h2b, 16'h4, 16'h6, 16'hfff8, 16'hfff6, 16'h16, 16'hffed, 16'h17, 16'h30, 16'h1b, 16'hffd5, 16'hffe7, 16'h89, 16'h6f, 16'hffdf, 16'hffda, 16'hffd6, 16'hffd7, 16'h63, 16'h74, 16'h23, 16'hffde, 16'hffdc, 16'h0, 16'hffa6, 16'hffdf, 16'h2c, 16'h45, 16'h34, 16'hffca, 16'hffab, 16'hffc0, 16'hb, 16'h4e, 16'h2b, 16'h17, 16'hffe8, 16'h1f, 16'h15, 16'h40, 16'h8, 16'h5, 16'hb, 16'hfff9, 16'hffef, 16'hff70, 16'hffa8, 16'hfff9, 16'hfffb, 16'h2b, 16'h3, 16'hff7a, 16'hff68, 16'hffe8, 16'hffd2, 16'hffd5, 16'hffe4, 16'hff80, 16'hff7e, 16'hfff8, 16'hfff9, 16'hffce, 16'hffd7, 16'hffd8, 16'hffd2, 16'h16, 16'h6, 16'hffdf, 16'hfffc, 16'h8, 16'h15, 16'h9, 16'h10, 16'h15, 16'h1d, 16'h10, 16'hf, 16'hfff9, 16'hff9c, 16'h55, 16'hbf, 16'had, 16'h54, 16'hffdf, 16'hffbc, 16'hffff, 16'h81, 16'h49, 16'hd, 16'h8, 16'he, 16'h10, 16'h1d, 16'h30, 16'h37, 16'hffd9, 16'hffd3, 16'h7, 16'hd, 16'h23, 16'h22, 16'hffd7, 16'hffaf, 16'hffb6, 16'hffed, 16'hffec, 16'h8, 16'hfffd, 16'hfff0, 16'hffbc, 16'hffa6, 16'hffd0, 16'hffe7, 16'hfff7, 16'h2, 16'h7, 16'hffcb, 16'hffff, 16'hfff1, 16'h19, 16'hfffd, 16'h44, 16'h8, 16'hffdf, 16'hfffa, 16'h8, 16'h35, 16'h37, 16'h7, 16'hfffd, 16'h0, 16'hffef, 16'h23, 16'h58, 16'h26, 16'hb, 16'hfffc, 16'hffee, 16'h3e, 16'h74, 16'h79, 16'h25, 16'h26, 16'h8, 16'h4, 16'h43, 16'h4f, 16'h44, 16'h41, 16'h1f, 16'ha, 16'h1c, 16'hffeb, 16'hffe9, 16'hffe0, 16'hfff6, 16'hffcd, 16'hfff5, 16'hffa2, 16'hffaf, 16'hffcb, 16'hffef, 16'hffe7, 16'hd, 16'hffcf, 16'hffdc, 16'hfff0, 16'h5c, 16'h43, 16'h60, 16'hfffe, 16'hb, 16'hf, 16'h46, 16'h51, 16'h47, 16'hffea, 16'hffee, 16'h5, 16'h1c, 16'h3b, 16'hfff7, 16'hffb9, 16'hffb0, 16'hffd1, 16'hffef, 16'hfffb, 16'hffef, 16'hfffb, 16'hffe3, 16'hffd3, 16'hfff7, 16'h19, 16'hffb1, 16'hffc0, 16'h1f, 16'hfffe, 16'hffef, 16'hffd9, 16'hffe8, 16'hffd4, 16'h6, 16'hffdf, 16'hffd5, 16'hffc8, 16'hffd6, 16'hfff5, 16'h19, 16'hffef, 16'hffef, 16'hffd8, 16'hffe0, 16'hfffe, 16'h15, 16'hffe6, 16'h4, 16'h4, 16'h16, 16'h12, 16'h16, 16'hfff4, 16'hffef, 16'hffa3, 16'hff8d, 16'h16, 16'h17, 16'hffc0, 16'hfffd, 16'hffb6, 16'hffd2, 16'h17, 16'hffef, 16'hffdf, 16'h23, 16'hffdf, 16'hfffa, 16'hb, 16'hfff1, 16'hffe1, 16'hffe9, 16'hffc5, 16'hfff0, 16'h16, 16'h1a, 16'hc, 16'h1, 16'hffdb, 16'h12, 16'hfff4, 16'hffef, 16'hffd8, 16'h1d, 16'hfffd, 16'hffe9, 16'hffbb, 16'hffd7, 16'hfffb, 16'h9, 16'hffd9, 16'h37, 16'h10, 16'hfff9, 16'h1, 16'h1, 16'hff83, 16'hff6b, 16'hffbe, 16'hffe0, 16'h1c, 16'hffdf, 16'hff77, 16'hff76, 16'hffb3, 16'hffd5, 16'h13, 16'hffe5, 16'hffd1, 16'hffc8, 16'hffe1, 16'h7, 16'h2b, 16'hffe8, 16'hffe1, 16'hffe4, 16'h11, 16'h1f, 16'h2c, 16'hfffa, 16'h1f, 16'h5, 16'h6, 16'h11, 16'h36, 16'h4, 16'hffe2, 16'hffd4, 16'hfffd, 16'hffca, 16'hffdc, 16'hfff1, 16'h4a, 16'h6, 16'hffae, 16'hffc7, 16'hffb2, 16'h16, 16'h64, 16'h58, 16'h9, 16'hffd4, 16'hffe1, 16'h23, 16'h84, 16'h80, 16'h38, 16'h9, 16'h1e, 16'h29, 16'h63, 16'h4a, 16'h22, 16'h11, 16'h16, 16'h21, 16'h25, 16'h8, 16'h8, 16'h31, 16'h21, 16'hfffe, 16'h3, 16'hffd4, 16'hffde, 16'hffa6, 16'hffc9, 16'hfffe, 16'h16, 16'hffa1, 16'hff8b, 16'hff4e, 16'hff53, 16'h33, 16'hffe1, 16'hffdc, 16'hffd4, 16'hffb3, 16'hffb1, 16'h3, 16'hffe3, 16'h0, 16'h17, 16'hc, 16'hffe7, 16'h17, 16'hfffb, 16'h43, 16'h51, 16'h34, 16'h33, 16'h10, 16'hffef, 16'h3a, 16'h3c, 16'h21, 16'h24, 16'h22, 16'h69, 16'hfff7, 16'hffa8, 16'hffec, 16'h30, 16'hffe9, 16'h28, 16'h1d, 16'hffec, 16'h31, 16'h42, 16'hffce, 16'hffdf, 16'hffc9, 16'hfff3, 16'h41, 16'h50, 16'hffa0, 16'hffc3, 16'hffaa, 16'hfff5, 16'hffdb, 16'hffc1, 16'hffc1, 16'hffb7, 16'hffba, 16'h12, 16'hffd9, 16'hffc3, 16'hffe0, 16'hffda, 16'h1d, 16'h2f, 16'hfffb, 16'hffbf, 16'h30, 16'h26, 16'hfff9, 16'h9, 16'h1b, 16'h33, 16'h11, 16'h2b, 16'hff8a, 16'hffbd, 16'h1, 16'hfff6, 16'h1f, 16'h4, 16'hfff4, 16'h2c, 16'h49, 16'hffff, 16'h3c, 16'hffe9, 16'h4a, 16'h5b, 16'h7d, 16'hffea, 16'h3f, 16'hffef, 16'h35, 16'h1b, 16'h20, 16'hfffa, 16'hfffa, 16'h23, 16'hffe6, 16'hffdf, 16'hffde, 16'hfff6, 16'h2a, 16'h7, 16'h6, 16'hfff7, 16'hffe3, 16'hfffc, 16'hfff8, 16'h1, 16'hffde, 16'hffe4, 16'hffc2, 16'hffe6, 16'hffd3, 16'hffc5, 16'hffbc, 16'hffd8, 16'hffc0, 16'hffc4, 16'hfffc, 16'hffe3, 16'hfff1, 16'hc, 16'hffea, 16'hffde, 16'hfff5, 16'h22, 16'h30, 16'h5c, 16'h1f, 16'hc, 16'h5, 16'h39, 16'h2e, 16'h80, 16'h3c, 16'h22, 16'hffce, 16'hffee, 16'h1c, 16'hffff, 16'hffca, 16'hfff5, 16'hffce, 16'hffe3, 16'h4e, 16'h4, 16'hfffb, 16'he, 16'hffce, 16'h8, 16'h5, 16'hffcc, 16'hffac, 16'hffdc, 16'hffce, 16'hffee, 16'hffcd, 16'hffb9, 16'hff9f, 16'h9, 16'hffe4, 16'hffd2, 16'hffe9, 16'hffcf, 16'hffdb, 16'hffd5, 16'hffca, 16'hffe3, 16'hffe2, 16'hffd4, 16'hffbd, 16'hffcf, 16'hfffe, 16'h5f, 16'h6b, 16'hffe6, 16'he, 16'hfffa, 16'h6, 16'h82, 16'h3b, 16'hfffc, 16'h28, 16'h24, 16'h8, 16'h4e, 16'h16, 16'hffe0, 16'hffe0, 16'hffc8, 16'hffe8, 16'hffe5, 16'hffc5, 16'hfff1, 16'hffe9, 16'hffc1, 16'hfff3, 16'hffd2, 16'hffc6, 16'hffe9, 16'h13, 16'hffdb, 16'hfffb, 16'hffe5, 16'h18, 16'h3b, 16'h3d, 16'h1a, 16'h34, 16'h51, 16'h19, 16'hfffe, 16'hfff4, 16'hfffe, 16'h12, 16'hc6, 16'hb9, 16'h66, 16'hffef, 16'he, 16'h14, 16'h61, 16'h63, 16'h1c, 16'hffe5, 16'hfffb, 16'hffc8, 16'hffdc, 16'hffcd, 16'hffb1, 16'hffcc, 16'hffc7, 16'hffd6, 16'hffd9, 16'hffca, 16'hffc8, 16'hffb4, 16'hffa6, 16'hffdd, 16'hfff4, 16'hffe6, 16'hffdc, 16'hffda, 16'hffbe, 16'hc, 16'hffed, 16'hffe2, 16'hffeb, 16'hffe2, 16'hfff2, 16'h6, 16'hff6c, 16'hffa5, 16'h45, 16'h1c, 16'h1a, 16'h3, 16'hff87, 16'hff91, 16'h22, 16'h0, 16'hffff, 16'h3, 16'hffa9, 16'hfff5, 16'hffd8, 16'hffcb, 16'hffb0, 16'h1e, 16'hffcd, 16'hfff9, 16'hffbe, 16'hffa6, 16'hffa0, 16'h11, 16'h5, 16'hfffa, 16'hff8d, 16'hff8e, 16'hff99, 16'hfffe, 16'he, 16'h10, 16'hffd4, 16'hffa5, 16'hffb2, 16'h20, 16'h0, 16'hffd8, 16'hff70, 16'hff71, 16'hff97, 16'h35, 16'h6, 16'hffcd, 16'hff8d, 16'hffa4, 16'hffa5, 16'h39, 16'hf, 16'hffd0, 16'hffbd, 16'hffdb, 16'hffdf, 16'h1b, 16'hffe7, 16'hff9a, 16'hff79, 16'hffb2, 16'hffee, 16'h2, 16'hfff6, 16'hffea, 16'hffb8, 16'hffef, 16'hfffe, 16'h2b, 16'h91, 16'h3a, 16'h2d, 16'h3a, 16'hffcc, 16'h1f, 16'h1a, 16'h59, 16'h51, 16'h18, 16'hffd8, 16'hffdc, 16'hffd9, 16'h22, 16'h2f, 16'h8, 16'h1, 16'h17, 16'hffee, 16'h1c, 16'h48, 16'h14, 16'h9, 16'h1d, 16'h14, 16'h1b, 16'h34, 16'hb, 16'hf, 16'h1d, 16'h30, 16'h2b, 16'h30, 16'h35, 16'ha, 16'hffd2, 16'hffb3, 16'h75, 16'h45, 16'h1c, 16'hffe8, 16'hffd4, 16'h18, 16'h74, 16'h58, 16'h52, 16'hffd9, 16'hffc2, 16'h24, 16'h7c, 16'h7d, 16'h8f, 16'h1a, 16'hffc8, 16'h28, 16'h7a, 16'h64, 16'h54, 16'hfffe, 16'hffd2, 16'h3f, 16'h69, 16'h4c, 16'ha, 16'hfffd, 16'hffa5, 16'hfffd, 16'h30, 16'h1e, 16'hfffb, 16'hffd3, 16'hffc5, 16'h1b, 16'hfff3, 16'hb, 16'hfffc, 16'h4, 16'h40, 16'h53, 16'h29, 16'h2, 16'hfff9, 16'hfff8, 16'h1, 16'h23, 16'h32, 16'hffe7, 16'hffea, 16'hfff4, 16'hffff, 16'hffee, 16'he, 16'hffcf, 16'hffd9, 16'hfff2, 16'h16, 16'h5, 16'h4, 16'hffe3, 16'hfff6, 16'h5, 16'hfff9, 16'hffff, 16'h6, 16'hfff9, 16'hffe4, 16'hffcd, 16'h4d, 16'h6, 16'hffcb, 16'h46, 16'h35, 16'h51, 16'h55, 16'hfff4, 16'h21, 16'h10, 16'hfffd, 16'h4e, 16'h24, 16'hfff2, 16'h28, 16'h12, 16'h21, 16'h4e, 16'h52, 16'hffd9, 16'hffec, 16'hfff0, 16'h2e, 16'h41, 16'h32, 16'h6, 16'hfffd, 16'h14, 16'h44, 16'h19, 16'h33, 16'h12, 16'h1e, 16'h26, 16'h17, 16'h23, 16'ha, 16'h2d, 16'h3f, 16'h2e, 16'h6, 16'h1, 16'hffd1, 16'hfff8, 16'h26, 16'h3b, 16'h6, 16'h2a, 16'hffd3, 16'hfff9, 16'h3b, 16'h2c, 16'h8, 16'ha, 16'hffde, 16'hffde, 16'hffff, 16'ha, 16'hf, 16'h29, 16'hffb9, 16'h2, 16'h6, 16'h13, 16'h3, 16'hd, 16'hffa8, 16'h10, 16'h31, 16'h34, 16'h17, 16'ha, 16'hffd8, 16'h9, 16'hffe6, 16'hffe0, 16'hfff2, 16'hffbc, 16'h2d, 16'h69, 16'h40, 16'hff9f, 16'hffa6, 16'hffb2, 16'hc, 16'h2, 16'h0, 16'hff7d, 16'hff9f, 16'hffc1, 16'hffec, 16'hff85, 16'hffb8, 16'hff99, 16'hffc6, 16'hffd0, 16'hfff7, 16'hffb6, 16'hffc9, 16'hffe8, 16'h15, 16'h1, 16'hfff2, 16'h3, 16'hfff1, 16'hfff5, 16'h5, 16'hfff9, 16'hffac, 16'h66, 16'haa, 16'h5c, 16'h5a, 16'hfff1, 16'hffc0, 16'h81, 16'hb4, 16'h61, 16'h2e, 16'he, 16'hffc8, 16'h3d, 16'h13, 16'h20, 16'h25, 16'h3b, 16'h4, 16'h65, 16'h41, 16'h2b, 16'h33, 16'h2c, 16'h12, 16'h72, 16'h3d, 16'h48, 16'h58, 16'h42, 16'hffe6, 16'h57, 16'h67, 16'h42, 16'h77, 16'h3, 16'hffa8, 16'hffb6, 16'h2b, 16'h40, 16'h1c, 16'h40, 16'hffe5, 16'hfffb, 16'h44, 16'h66, 16'h1f, 16'h1c, 16'hffd0, 16'hffce, 16'h25, 16'h45, 16'h32, 16'h20, 16'hffaf, 16'h2, 16'h1f, 16'h3d, 16'h30, 16'h6, 16'hffeb, 16'hffcf, 16'hfff4, 16'h37, 16'h37, 16'h36, 16'hffd1, 16'hffcf, 16'h1c, 16'h2d, 16'h45, 16'h23, 16'hffe3, 16'hffe0, 16'hffe5, 16'hffe7, 16'hffd6, 16'hffcd, 16'h31, 16'h3d, 16'h37, 16'h4, 16'hffdf, 16'hffb9, 16'h0, 16'h1b, 16'h18, 16'hffe5, 16'hff90, 16'hff7c, 16'hffc8, 16'hffac, 16'hff79, 16'hffab, 16'hff78, 16'hff92, 16'hffad, 16'hff88, 16'hff92, 16'hffec, 16'hffd8, 16'hffef, 16'h8, 16'hffdf, 16'h1d, 16'h68, 16'h58, 16'h33, 16'hffd9, 16'hffe4, 16'h17, 16'h57, 16'h60, 16'h10, 16'hffdf, 16'hfff7, 16'hfff3, 16'h38, 16'h5d, 16'h24, 16'h7, 16'h24, 16'h23, 16'h50, 16'h58, 16'h44, 16'hffd5, 16'h6, 16'h58, 16'h48, 16'h4e, 16'h17, 16'h11, 16'hfff2, 16'h2, 16'hffdd, 16'hffb1, 16'h1, 16'hffff, 16'hffe9, 16'hfff0, 16'hffab, 16'hffb4, 16'hfff2, 16'h1, 16'hffee, 16'hffbf, 16'hffc2, 16'hffe9, 16'hc, 16'hffd9, 16'h11, 16'h2, 16'hffe6, 16'h2f, 16'h24, 16'h35, 16'h4c, 16'h25, 16'h28, 16'ha, 16'h2, 16'h30, 16'hffff, 16'hffdb, 16'hffff, 16'h27, 16'h12, 16'hffd9, 16'hffd1, 16'hffdd, 16'h1e, 16'h56, 16'h15, 16'hffe6, 16'hffbe, 16'ha, 16'h76, 16'h95, 16'hf, 16'h4, 16'h27, 16'hffe1, 16'hffdb, 16'hfffc, 16'h14, 16'h21, 16'hffe1, 16'hfff7, 16'h13, 16'h13, 16'hfff4, 16'h2b, 16'hffd0, 16'hf, 16'h16, 16'h0, 16'h1a, 16'hffeb, 16'h29, 16'h4e, 16'h1, 16'h0, 16'h18, 16'hffeb, 16'hfffb, 16'h1a, 16'hfff6, 16'h6, 16'h22, 16'h27, 16'hd, 16'h19, 16'hfff9, 16'h14, 16'h17, 16'h3, 16'hffd7, 16'h9, 16'h20, 16'h18, 16'h12, 16'h26, 16'h1e, 16'h30, 16'hc, 16'hc, 16'h5, 16'hffde, 16'hffe2, 16'h2b, 16'h9, 16'h1, 16'hffea, 16'hfff3, 16'hffe0, 16'hffc5, 16'hfff8, 16'h5, 16'ha, 16'hffdb, 16'hffdd, 16'hffad, 16'hffec, 16'hf, 16'h40, 16'hffe5, 16'hffda, 16'hfff5, 16'h5a, 16'h53, 16'h56, 16'hffea, 16'hffe6, 16'h4, 16'hfff3, 16'h22, 16'hd, 16'hffef, 16'hffb2, 16'hffcf, 16'hfff4, 16'h8, 16'h0, 16'h5, 16'h2, 16'h2, 16'hffe2, 16'hffe0, 16'hffc2, 16'hffe7, 16'hfffd, 16'h7, 16'hffd7, 16'hffe4, 16'hffd1, 16'hffe5, 16'hffde, 16'hfff6, 16'hffef, 16'hb, 16'h12, 16'hffcc, 16'hffb3, 16'hfffb, 16'hffd9, 16'hc, 16'h28, 16'h12, 16'hfff5, 16'h33, 16'h3b, 16'h6c, 16'hfff8, 16'h14, 16'h3b, 16'h92, 16'h86, 16'h3b, 16'h27, 16'hfffd, 16'h69, 16'h4f, 16'h11, 16'hffe6, 16'h4, 16'hfff2, 16'hfffd, 16'hfff2, 16'hfff3, 16'hfff0, 16'hd, 16'h8, 16'hffc7, 16'hfff1, 16'hffe4, 16'hffdf, 16'hffea, 16'hffd1, 16'hffde, 16'h3, 16'hffca, 16'hffb5, 16'hffee, 16'hffed, 16'hfffc, 16'h9, 16'h0, 16'h2e, 16'h5a, 16'hffec, 16'hffdc, 16'h24, 16'h3b, 16'h5d, 16'h76, 16'h10, 16'hffd6, 16'h46, 16'h40, 16'h3e, 16'h60, 16'h6, 16'hfff2, 16'h31, 16'h37, 16'h4c, 16'h56, 16'hfff2, 16'hfff4, 16'hffae, 16'hffc4, 16'hffd8, 16'h4f, 16'hffe0, 16'hc, 16'hffd7, 16'hffa9, 16'hffe9, 16'h41};
    // logic signed [15:0] threshold [0:OC-1] = {-16'd31, -16'd73, -16'd16, -16'd33, -16'd13, -16'd3, -16'd1543, -16'd4, -16'd8, -16'd14};
    logic [CONV1_IMG_OUT_SIZE*CONV1_IMG_OUT_SIZE-1:0] conv1_img_out [0:CONV1_OC-1];
    logic [POOL1_IMG_OUT_SIZE*POOL1_IMG_OUT_SIZE-1:0] pool1_img_out [0:CONV1_OC-1];
    logic [CONV2_IMG_OUT_SIZE*CONV2_IMG_OUT_SIZE-1:0] conv2_img_out [0:CONV2_OC-1];
    logic [POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE-1:0] pool2_img_out [0:CONV2_OC-1];
    logic [FC_IC-1:0] fc_in;
    logic signed [15:0] fc_out [0:FC_OC-1];
    logic conv1_data_ready;
    logic pool1_data_ready;
    logic conv2_data_ready;
    logic pool2_data_ready;
    logic fc_data_ready;

    Conv2d #(
        .IC(CONV1_IC),
        .OC(CONV1_OC),
        .IMG_IN_SIZE(CONV1_IMG_IN_SIZE)
    ) conv1 (
        .clk(clk),
        .data_in_ready(data_in_ready),
        .img_in(conv1_img_in),
        .weights(conv1_weights),
        .img_out(conv1_img_out),
        .data_out_ready(conv1_data_ready)
    );

    MaxPool2d #(
        .IC(CONV1_OC),
        .IMG_IN_SIZE(CONV1_IMG_OUT_SIZE)
    ) pool1 (
        .clk(clk),
        .data_in_ready(conv1_data_ready),
        .img_in(conv1_img_out),
        .img_out(pool1_img_out),
        .data_out_ready(pool1_data_ready)
    );

    Conv2d #(
        .IC(CONV1_OC),
        .OC(CONV2_OC),
        .IMG_IN_SIZE(POOL1_IMG_OUT_SIZE)
    ) conv2 (
        .clk(clk),
        .data_in_ready(pool1_data_ready),
        .img_in(pool1_img_out),
        .weights(conv2_weights),
        .img_out(conv2_img_out),
        .data_out_ready(conv2_data_ready)
    );

    MaxPool2d #(
        .IC(CONV2_OC),
        .IMG_IN_SIZE(CONV2_IMG_OUT_SIZE)
    ) pool2 (
        .clk(clk),
        .data_in_ready(conv2_data_ready),
        .img_in(conv2_img_out),
        .img_out(pool2_img_out),
        .data_out_ready(pool2_data_ready)
    );

    genvar conv2_oc;
    generate
        for (conv2_oc=0; conv2_oc<CONV2_OC; conv2_oc=conv2_oc+1) begin
            assign fc_in[conv2_oc*POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE +: POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE] = pool2_img_out[conv2_oc];
        end
    endgenerate

    FC #(
        .IC(FC_IC),
        .OC(FC_OC)
    ) fc (
        .clk(clk),
        .data_in_ready(pool2_data_ready),
        .in(fc_in),
        .weights(fc_weights),
        .out(fc_out),
        .data_out_ready(fc_data_ready)
    );

    Comparator #(
        .IC(FC_OC),
    ) compare (
        .clk(clk),
        .data_in_ready(fc_data_ready),
        .in(fc_out),
        .out(result),
        .data_out_ready(data_out_ready)
    );

    // wire _unused_ok = &{result};

endmodule

